module odo_apply_pbox1(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[6] = in[0];
    assign out[484] = in[1];
    assign out[367] = in[2];
    assign out[347] = in[3];
    assign out[69] = in[4];
    assign out[597] = in[5];
    assign out[68] = in[6];
    assign out[112] = in[7];
    assign out[73] = in[8];
    assign out[380] = in[9];
    assign out[429] = in[10];
    assign out[508] = in[11];
    assign out[140] = in[12];
    assign out[296] = in[13];
    assign out[617] = in[14];
    assign out[458] = in[15];
    assign out[385] = in[16];
    assign out[130] = in[17];
    assign out[384] = in[18];
    assign out[547] = in[19];
    assign out[613] = in[20];
    assign out[185] = in[21];
    assign out[604] = in[22];
    assign out[266] = in[23];
    assign out[467] = in[24];
    assign out[2] = in[25];
    assign out[57] = in[26];
    assign out[4] = in[27];
    assign out[407] = in[28];
    assign out[99] = in[29];
    assign out[193] = in[30];
    assign out[144] = in[31];
    assign out[550] = in[32];
    assign out[31] = in[33];
    assign out[104] = in[34];
    assign out[33] = in[35];
    assign out[565] = in[36];
    assign out[280] = in[37];
    assign out[526] = in[38];
    assign out[340] = in[39];
    assign out[343] = in[40];
    assign out[486] = in[41];
    assign out[43] = in[42];
    assign out[235] = in[43];
    assign out[324] = in[44];
    assign out[348] = in[45];
    assign out[283] = in[46];
    assign out[466] = in[47];
    assign out[417] = in[48];
    assign out[428] = in[49];
    assign out[238] = in[50];
    assign out[164] = in[51];
    assign out[631] = in[52];
    assign out[54] = in[53];
    assign out[153] = in[54];
    assign out[410] = in[55];
    assign out[638] = in[56];
    assign out[24] = in[57];
    assign out[113] = in[58];
    assign out[302] = in[59];
    assign out[361] = in[60];
    assign out[28] = in[61];
    assign out[29] = in[62];
    assign out[247] = in[63];
    assign out[445] = in[64];
    assign out[56] = in[65];
    assign out[485] = in[66];
    assign out[446] = in[67];
    assign out[498] = in[68];
    assign out[488] = in[69];
    assign out[371] = in[70];
    assign out[308] = in[71];
    assign out[600] = in[72];
    assign out[255] = in[73];
    assign out[602] = in[74];
    assign out[494] = in[75];
    assign out[530] = in[76];
    assign out[394] = in[77];
    assign out[529] = in[78];
    assign out[199] = in[79];
    assign out[204] = in[80];
    assign out[260] = in[81];
    assign out[533] = in[82];
    assign out[262] = in[83];
    assign out[125] = in[84];
    assign out[83] = in[85];
    assign out[401] = in[86];
    assign out[64] = in[87];
    assign out[542] = in[88];
    assign out[513] = in[89];
    assign out[3] = in[90];
    assign out[190] = in[91];
    assign out[473] = in[92];
    assign out[448] = in[93];
    assign out[409] = in[94];
    assign out[155] = in[95];
    assign out[475] = in[96];
    assign out[561] = in[97];
    assign out[197] = in[98];
    assign out[628] = in[99];
    assign out[551] = in[100];
    assign out[320] = in[101];
    assign out[326] = in[102];
    assign out[420] = in[103];
    assign out[46] = in[104];
    assign out[82] = in[105];
    assign out[142] = in[106];
    assign out[108] = in[107];
    assign out[236] = in[108];
    assign out[333] = in[109];
    assign out[44] = in[110];
    assign out[160] = in[111];
    assign out[470] = in[112];
    assign out[114] = in[113];
    assign out[287] = in[114];
    assign out[432] = in[115];
    assign out[107] = in[116];
    assign out[171] = in[117];
    assign out[154] = in[118];
    assign out[168] = in[119];
    assign out[344] = in[120];
    assign out[358] = in[121];
    assign out[221] = in[122];
    assign out[36] = in[123];
    assign out[58] = in[124];
    assign out[440] = in[125];
    assign out[492] = in[126];
    assign out[591] = in[127];
    assign out[227] = in[128];
    assign out[393] = in[129];
    assign out[129] = in[130];
    assign out[161] = in[131];
    assign out[345] = in[132];
    assign out[584] = in[133];
    assign out[517] = in[134];
    assign out[399] = in[135];
    assign out[523] = in[136];
    assign out[489] = in[137];
    assign out[522] = in[138];
    assign out[559] = in[139];
    assign out[605] = in[140];
    assign out[323] = in[141];
    assign out[120] = in[142];
    assign out[594] = in[143];
    assign out[609] = in[144];
    assign out[241] = in[145];
    assign out[49] = in[146];
    assign out[400] = in[147];
    assign out[126] = in[148];
    assign out[285] = in[149];
    assign out[570] = in[150];
    assign out[538] = in[151];
    assign out[603] = in[152];
    assign out[537] = in[153];
    assign out[354] = in[154];
    assign out[65] = in[155];
    assign out[305] = in[156];
    assign out[474] = in[157];
    assign out[500] = in[158];
    assign out[546] = in[159];
    assign out[200] = in[160];
    assign out[544] = in[161];
    assign out[311] = in[162];
    assign out[17] = in[163];
    assign out[481] = in[164];
    assign out[184] = in[165];
    assign out[80] = in[166];
    assign out[303] = in[167];
    assign out[555] = in[168];
    assign out[18] = in[169];
    assign out[624] = in[170];
    assign out[201] = in[171];
    assign out[637] = in[172];
    assign out[464] = in[173];
    assign out[209] = in[174];
    assign out[141] = in[175];
    assign out[378] = in[176];
    assign out[437] = in[177];
    assign out[438] = in[178];
    assign out[535] = in[179];
    assign out[220] = in[180];
    assign out[136] = in[181];
    assign out[636] = in[182];
    assign out[365] = in[183];
    assign out[472] = in[184];
    assign out[449] = in[185];
    assign out[587] = in[186];
    assign out[574] = in[187];
    assign out[363] = in[188];
    assign out[480] = in[189];
    assign out[450] = in[190];
    assign out[592] = in[191];
    assign out[639] = in[192];
    assign out[169] = in[193];
    assign out[520] = in[194];
    assign out[150] = in[195];
    assign out[579] = in[196];
    assign out[580] = in[197];
    assign out[47] = in[198];
    assign out[589] = in[199];
    assign out[583] = in[200];
    assign out[273] = in[201];
    assign out[416] = in[202];
    assign out[42] = in[203];
    assign out[418] = in[204];
    assign out[496] = in[205];
    assign out[355] = in[206];
    assign out[117] = in[207];
    assign out[499] = in[208];
    assign out[249] = in[209];
    assign out[593] = in[210];
    assign out[121] = in[211];
    assign out[426] = in[212];
    assign out[232] = in[213];
    assign out[63] = in[214];
    assign out[598] = in[215];
    assign out[290] = in[216];
    assign out[540] = in[217];
    assign out[173] = in[218];
    assign out[330] = in[219];
    assign out[539] = in[220];
    assign out[295] = in[221];
    assign out[482] = in[222];
    assign out[191] = in[223];
    assign out[282] = in[224];
    assign out[548] = in[225];
    assign out[364] = in[226];
    assign out[519] = in[227];
    assign out[286] = in[228];
    assign out[276] = in[229];
    assign out[366] = in[230];
    assign out[77] = in[231];
    assign out[633] = in[232];
    assign out[457] = in[233];
    assign out[288] = in[234];
    assign out[139] = in[235];
    assign out[425] = in[236];
    assign out[497] = in[237];
    assign out[502] = in[238];
    assign out[207] = in[239];
    assign out[312] = in[240];
    assign out[352] = in[241];
    assign out[91] = in[242];
    assign out[379] = in[243];
    assign out[243] = in[244];
    assign out[211] = in[245];
    assign out[32] = in[246];
    assign out[332] = in[247];
    assign out[462] = in[248];
    assign out[270] = in[249];
    assign out[413] = in[250];
    assign out[219] = in[251];
    assign out[388] = in[252];
    assign out[545] = in[253];
    assign out[225] = in[254];
    assign out[405] = in[255];
    assign out[179] = in[256];
    assign out[230] = in[257];
    assign out[532] = in[258];
    assign out[127] = in[259];
    assign out[251] = in[260];
    assign out[325] = in[261];
    assign out[189] = in[262];
    assign out[611] = in[263];
    assign out[186] = in[264];
    assign out[252] = in[265];
    assign out[614] = in[266];
    assign out[477] = in[267];
    assign out[493] = in[268];
    assign out[119] = in[269];
    assign out[192] = in[270];
    assign out[618] = in[271];
    assign out[291] = in[272];
    assign out[131] = in[273];
    assign out[629] = in[274];
    assign out[76] = in[275];
    assign out[373] = in[276];
    assign out[341] = in[277];
    assign out[375] = in[278];
    assign out[19] = in[279];
    assign out[143] = in[280];
    assign out[208] = in[281];
    assign out[406] = in[282];
    assign out[521] = in[283];
    assign out[165] = in[284];
    assign out[377] = in[285];
    assign out[23] = in[286];
    assign out[315] = in[287];
    assign out[571] = in[288];
    assign out[216] = in[289];
    assign out[105] = in[290];
    assign out[501] = in[291];
    assign out[215] = in[292];
    assign out[93] = in[293];
    assign out[567] = in[294];
    assign out[632] = in[295];
    assign out[278] = in[296];
    assign out[588] = in[297];
    assign out[444] = in[298];
    assign out[573] = in[299];
    assign out[145] = in[300];
    assign out[87] = in[301];
    assign out[585] = in[302];
    assign out[118] = in[303];
    assign out[304] = in[304];
    assign out[543] = in[305];
    assign out[608] = in[306];
    assign out[495] = in[307];
    assign out[40] = in[308];
    assign out[182] = in[309];
    assign out[356] = in[310];
    assign out[453] = in[311];
    assign out[157] = in[312];
    assign out[424] = in[313];
    assign out[187] = in[314];
    assign out[51] = in[315];
    assign out[256] = in[316];
    assign out[226] = in[317];
    assign out[5] = in[318];
    assign out[461] = in[319];
    assign out[7] = in[320];
    assign out[612] = in[321];
    assign out[549] = in[322];
    assign out[59] = in[323];
    assign out[626] = in[324];
    assign out[439] = in[325];
    assign out[536] = in[326];
    assign out[610] = in[327];
    assign out[374] = in[328];
    assign out[202] = in[329];
    assign out[67] = in[330];
    assign out[541] = in[331];
    assign out[507] = in[332];
    assign out[430] = in[333];
    assign out[338] = in[334];
    assign out[86] = in[335];
    assign out[135] = in[336];
    assign out[196] = in[337];
    assign out[307] = in[338];
    assign out[386] = in[339];
    assign out[203] = in[340];
    assign out[250] = in[341];
    assign out[516] = in[342];
    assign out[1] = in[343];
    assign out[518] = in[344];
    assign out[564] = in[345];
    assign out[346] = in[346];
    assign out[205] = in[347];
    assign out[84] = in[348];
    assign out[576] = in[349];
    assign out[319] = in[350];
    assign out[578] = in[351];
    assign out[321] = in[352];
    assign out[562] = in[353];
    assign out[217] = in[354];
    assign out[337] = in[355];
    assign out[229] = in[356];
    assign out[293] = in[357];
    assign out[34] = in[358];
    assign out[27] = in[359];
    assign out[300] = in[360];
    assign out[224] = in[361];
    assign out[98] = in[362];
    assign out[95] = in[363];
    assign out[163] = in[364];
    assign out[369] = in[365];
    assign out[490] = in[366];
    assign out[322] = in[367];
    assign out[149] = in[368];
    assign out[515] = in[369];
    assign out[590] = in[370];
    assign out[389] = in[371];
    assign out[166] = in[372];
    assign out[172] = in[373];
    assign out[471] = in[374];
    assign out[97] = in[375];
    assign out[239] = in[376];
    assign out[268] = in[377];
    assign out[237] = in[378];
    assign out[178] = in[379];
    assign out[38] = in[380];
    assign out[272] = in[381];
    assign out[55] = in[382];
    assign out[228] = in[383];
    assign out[625] = in[384];
    assign out[188] = in[385];
    assign out[147] = in[386];
    assign out[12] = in[387];
    assign out[505] = in[388];
    assign out[566] = in[389];
    assign out[621] = in[390];
    assign out[101] = in[391];
    assign out[569] = in[392];
    assign out[218] = in[393];
    assign out[524] = in[394];
    assign out[20] = in[395];
    assign out[382] = in[396];
    assign out[478] = in[397];
    assign out[11] = in[398];
    assign out[257] = in[399];
    assign out[110] = in[400];
    assign out[514] = in[401];
    assign out[455] = in[402];
    assign out[318] = in[403];
    assign out[132] = in[404];
    assign out[21] = in[405];
    assign out[45] = in[406];
    assign out[601] = in[407];
    assign out[404] = in[408];
    assign out[510] = in[409];
    assign out[586] = in[410];
    assign out[88] = in[411];
    assign out[89] = in[412];
    assign out[148] = in[413];
    assign out[213] = in[414];
    assign out[240] = in[415];
    assign out[469] = in[416];
    assign out[328] = in[417];
    assign out[615] = in[418];
    assign out[158] = in[419];
    assign out[267] = in[420];
    assign out[534] = in[421];
    assign out[269] = in[422];
    assign out[572] = in[423];
    assign out[223] = in[424];
    assign out[41] = in[425];
    assign out[284] = in[426];
    assign out[70] = in[427];
    assign out[398] = in[428];
    assign out[463] = in[429];
    assign out[281] = in[430];
    assign out[607] = in[431];
    assign out[231] = in[432];
    assign out[563] = in[433];
    assign out[90] = in[434];
    assign out[81] = in[435];
    assign out[331] = in[436];
    assign out[134] = in[437];
    assign out[292] = in[438];
    assign out[174] = in[439];
    assign out[362] = in[440];
    assign out[554] = in[441];
    assign out[122] = in[442];
    assign out[242] = in[443];
    assign out[100] = in[444];
    assign out[575] = in[445];
    assign out[483] = in[446];
    assign out[342] = in[447];
    assign out[94] = in[448];
    assign out[210] = in[449];
    assign out[423] = in[450];
    assign out[309] = in[451];
    assign out[306] = in[452];
    assign out[35] = in[453];
    assign out[15] = in[454];
    assign out[183] = in[455];
    assign out[8] = in[456];
    assign out[103] = in[457];
    assign out[451] = in[458];
    assign out[381] = in[459];
    assign out[263] = in[460];
    assign out[13] = in[461];
    assign out[37] = in[462];
    assign out[314] = in[463];
    assign out[212] = in[464];
    assign out[397] = in[465];
    assign out[244] = in[466];
    assign out[298] = in[467];
    assign out[60] = in[468];
    assign out[133] = in[469];
    assign out[248] = in[470];
    assign out[206] = in[471];
    assign out[115] = in[472];
    assign out[116] = in[473];
    assign out[264] = in[474];
    assign out[50] = in[475];
    assign out[279] = in[476];
    assign out[52] = in[477];
    assign out[265] = in[478];
    assign out[310] = in[479];
    assign out[334] = in[480];
    assign out[30] = in[481];
    assign out[411] = in[482];
    assign out[350] = in[483];
    assign out[390] = in[484];
    assign out[316] = in[485];
    assign out[78] = in[486];
    assign out[277] = in[487];
    assign out[335] = in[488];
    assign out[619] = in[489];
    assign out[479] = in[490];
    assign out[557] = in[491];
    assign out[622] = in[492];
    assign out[606] = in[493];
    assign out[261] = in[494];
    assign out[427] = in[495];
    assign out[75] = in[496];
    assign out[630] = in[497];
    assign out[246] = in[498];
    assign out[74] = in[499];
    assign out[351] = in[500];
    assign out[53] = in[501];
    assign out[431] = in[502];
    assign out[392] = in[503];
    assign out[525] = in[504];
    assign out[180] = in[505];
    assign out[435] = in[506];
    assign out[396] = in[507];
    assign out[128] = in[508];
    assign out[376] = in[509];
    assign out[25] = in[510];
    assign out[436] = in[511];
    assign out[422] = in[512];
    assign out[123] = in[513];
    assign out[558] = in[514];
    assign out[476] = in[515];
    assign out[175] = in[516];
    assign out[349] = in[517];
    assign out[454] = in[518];
    assign out[62] = in[519];
    assign out[468] = in[520];
    assign out[0] = in[521];
    assign out[124] = in[522];
    assign out[329] = in[523];
    assign out[568] = in[524];
    assign out[531] = in[525];
    assign out[48] = in[526];
    assign out[176] = in[527];
    assign out[289] = in[528];
    assign out[465] = in[529];
    assign out[336] = in[530];
    assign out[620] = in[531];
    assign out[274] = in[532];
    assign out[156] = in[533];
    assign out[66] = in[534];
    assign out[253] = in[535];
    assign out[9] = in[536];
    assign out[447] = in[537];
    assign out[357] = in[538];
    assign out[61] = in[539];
    assign out[22] = in[540];
    assign out[146] = in[541];
    assign out[85] = in[542];
    assign out[491] = in[543];
    assign out[553] = in[544];
    assign out[433] = in[545];
    assign out[151] = in[546];
    assign out[353] = in[547];
    assign out[528] = in[548];
    assign out[198] = in[549];
    assign out[511] = in[550];
    assign out[275] = in[551];
    assign out[10] = in[552];
    assign out[138] = in[553];
    assign out[560] = in[554];
    assign out[301] = in[555];
    assign out[317] = in[556];
    assign out[222] = in[557];
    assign out[245] = in[558];
    assign out[102] = in[559];
    assign out[39] = in[560];
    assign out[634] = in[561];
    assign out[259] = in[562];
    assign out[460] = in[563];
    assign out[233] = in[564];
    assign out[635] = in[565];
    assign out[599] = in[566];
    assign out[254] = in[567];
    assign out[26] = in[568];
    assign out[106] = in[569];
    assign out[595] = in[570];
    assign out[577] = in[571];
    assign out[195] = in[572];
    assign out[111] = in[573];
    assign out[271] = in[574];
    assign out[459] = in[575];
    assign out[556] = in[576];
    assign out[487] = in[577];
    assign out[372] = in[578];
    assign out[403] = in[579];
    assign out[258] = in[580];
    assign out[327] = in[581];
    assign out[370] = in[582];
    assign out[313] = in[583];
    assign out[339] = in[584];
    assign out[527] = in[585];
    assign out[181] = in[586];
    assign out[395] = in[587];
    assign out[421] = in[588];
    assign out[71] = in[589];
    assign out[414] = in[590];
    assign out[616] = in[591];
    assign out[177] = in[592];
    assign out[72] = in[593];
    assign out[402] = in[594];
    assign out[299] = in[595];
    assign out[442] = in[596];
    assign out[443] = in[597];
    assign out[623] = in[598];
    assign out[360] = in[599];
    assign out[503] = in[600];
    assign out[581] = in[601];
    assign out[441] = in[602];
    assign out[506] = in[603];
    assign out[359] = in[604];
    assign out[387] = in[605];
    assign out[137] = in[606];
    assign out[415] = in[607];
    assign out[167] = in[608];
    assign out[194] = in[609];
    assign out[552] = in[610];
    assign out[79] = in[611];
    assign out[16] = in[612];
    assign out[582] = in[613];
    assign out[434] = in[614];
    assign out[383] = in[615];
    assign out[504] = in[616];
    assign out[96] = in[617];
    assign out[159] = in[618];
    assign out[92] = in[619];
    assign out[14] = in[620];
    assign out[627] = in[621];
    assign out[391] = in[622];
    assign out[456] = in[623];
    assign out[214] = in[624];
    assign out[509] = in[625];
    assign out[152] = in[626];
    assign out[596] = in[627];
    assign out[294] = in[628];
    assign out[170] = in[629];
    assign out[412] = in[630];
    assign out[297] = in[631];
    assign out[452] = in[632];
    assign out[234] = in[633];
    assign out[512] = in[634];
    assign out[109] = in[635];
    assign out[162] = in[636];
    assign out[419] = in[637];
    assign out[368] = in[638];
    assign out[408] = in[639];
endmodule

