module odo_encrypt_loop(clk, in, read, out, write);
    input clk;
    input [639:0] in;
    input read;
    output reg [639:0] out;
    output write;
    reg [639:0] state[9:0];
    wire [639:0] next[9:0];
    always @(posedge clk) state[1] <= next[0];
    always @(posedge clk) state[2] <= next[1];
    always @(posedge clk) state[3] <= next[2];
    always @(posedge clk) state[4] <= next[3];
    always @(posedge clk) state[5] <= next[4];
    always @(posedge clk) state[6] <= next[5];
    always @(posedge clk) state[7] <= next[6];
    always @(posedge clk) state[8] <= next[7];
    always @(posedge clk) state[9] <= next[8];
    assign next[9] = state[9];
    wire [9:0] roundkey[8:0];
    reg [3:0] period[18:0];
    always @(posedge clk) period[1] <= period[0];
    always @(posedge clk) period[2] <= period[1];
    always @(posedge clk) period[3] <= period[2];
    always @(posedge clk) period[4] <= period[3];
    always @(posedge clk) period[5] <= period[4];
    always @(posedge clk) period[6] <= period[5];
    always @(posedge clk) period[7] <= period[6];
    always @(posedge clk) period[8] <= period[7];
    always @(posedge clk) period[9] <= period[8];
    always @(posedge clk) period[10] <= period[9];
    always @(posedge clk) period[11] <= period[10];
    always @(posedge clk) period[12] <= period[11];
    always @(posedge clk) period[13] <= period[12];
    always @(posedge clk) period[14] <= period[13];
    always @(posedge clk) period[15] <= period[14];
    always @(posedge clk) period[16] <= period[15];
    always @(posedge clk) period[17] <= period[16];
    always @(posedge clk) period[18] <= period[17];
    odo_get_round_key0 get_key0(clk, period[0], roundkey[0]);
    odo_full_round round0(clk, roundkey[0], state[0], next[0]);
    odo_get_round_key1 get_key1(clk, period[2], roundkey[1]);
    odo_full_round round1(clk, roundkey[1], state[1], next[1]);
    odo_get_round_key2 get_key2(clk, period[4], roundkey[2]);
    odo_full_round round2(clk, roundkey[2], state[2], next[2]);
    odo_get_round_key3 get_key3(clk, period[6], roundkey[3]);
    odo_full_round round3(clk, roundkey[3], state[3], next[3]);
    odo_get_round_key4 get_key4(clk, period[8], roundkey[4]);
    odo_full_round round4(clk, roundkey[4], state[4], next[4]);
    odo_get_round_key5 get_key5(clk, period[10], roundkey[5]);
    odo_full_round round5(clk, roundkey[5], state[5], next[5]);
    odo_get_round_key6 get_key6(clk, period[12], roundkey[6]);
    odo_full_round round6(clk, roundkey[6], state[6], next[6]);
    odo_get_round_key7 get_key7(clk, period[14], roundkey[7]);
    odo_full_round round7(clk, roundkey[7], state[7], next[7]);
    odo_get_round_key8 get_key8(clk, period[16], roundkey[8]);
    odo_full_round round8(clk, roundkey[8], state[8], next[8]);
    always @(posedge clk) begin
        if (read)
        begin
            period[0] <= 0;
            state[0] <= in;
        end
        else
        begin
            period[0] <= period[18]+1;
            state[0] <= next[9];
        end
        out <= next[2];
    end
    reg [177:0] progress;
    initial progress = 178'h0;
    always @(posedge clk) progress[0] <= read;
    always @(posedge clk) progress[1] <= progress[0];
    always @(posedge clk) progress[2] <= progress[1];
    always @(posedge clk) progress[3] <= progress[2];
    always @(posedge clk) progress[4] <= progress[3];
    always @(posedge clk) progress[5] <= progress[4];
    always @(posedge clk) progress[6] <= progress[5];
    always @(posedge clk) progress[7] <= progress[6];
    always @(posedge clk) progress[8] <= progress[7];
    always @(posedge clk) progress[9] <= progress[8];
    always @(posedge clk) progress[10] <= progress[9];
    always @(posedge clk) progress[11] <= progress[10];
    always @(posedge clk) progress[12] <= progress[11];
    always @(posedge clk) progress[13] <= progress[12];
    always @(posedge clk) progress[14] <= progress[13];
    always @(posedge clk) progress[15] <= progress[14];
    always @(posedge clk) progress[16] <= progress[15];
    always @(posedge clk) progress[17] <= progress[16];
    always @(posedge clk) progress[18] <= progress[17];
    always @(posedge clk) progress[19] <= progress[18];
    always @(posedge clk) progress[20] <= progress[19];
    always @(posedge clk) progress[21] <= progress[20];
    always @(posedge clk) progress[22] <= progress[21];
    always @(posedge clk) progress[23] <= progress[22];
    always @(posedge clk) progress[24] <= progress[23];
    always @(posedge clk) progress[25] <= progress[24];
    always @(posedge clk) progress[26] <= progress[25];
    always @(posedge clk) progress[27] <= progress[26];
    always @(posedge clk) progress[28] <= progress[27];
    always @(posedge clk) progress[29] <= progress[28];
    always @(posedge clk) progress[30] <= progress[29];
    always @(posedge clk) progress[31] <= progress[30];
    always @(posedge clk) progress[32] <= progress[31];
    always @(posedge clk) progress[33] <= progress[32];
    always @(posedge clk) progress[34] <= progress[33];
    always @(posedge clk) progress[35] <= progress[34];
    always @(posedge clk) progress[36] <= progress[35];
    always @(posedge clk) progress[37] <= progress[36];
    always @(posedge clk) progress[38] <= progress[37];
    always @(posedge clk) progress[39] <= progress[38];
    always @(posedge clk) progress[40] <= progress[39];
    always @(posedge clk) progress[41] <= progress[40];
    always @(posedge clk) progress[42] <= progress[41];
    always @(posedge clk) progress[43] <= progress[42];
    always @(posedge clk) progress[44] <= progress[43];
    always @(posedge clk) progress[45] <= progress[44];
    always @(posedge clk) progress[46] <= progress[45];
    always @(posedge clk) progress[47] <= progress[46];
    always @(posedge clk) progress[48] <= progress[47];
    always @(posedge clk) progress[49] <= progress[48];
    always @(posedge clk) progress[50] <= progress[49];
    always @(posedge clk) progress[51] <= progress[50];
    always @(posedge clk) progress[52] <= progress[51];
    always @(posedge clk) progress[53] <= progress[52];
    always @(posedge clk) progress[54] <= progress[53];
    always @(posedge clk) progress[55] <= progress[54];
    always @(posedge clk) progress[56] <= progress[55];
    always @(posedge clk) progress[57] <= progress[56];
    always @(posedge clk) progress[58] <= progress[57];
    always @(posedge clk) progress[59] <= progress[58];
    always @(posedge clk) progress[60] <= progress[59];
    always @(posedge clk) progress[61] <= progress[60];
    always @(posedge clk) progress[62] <= progress[61];
    always @(posedge clk) progress[63] <= progress[62];
    always @(posedge clk) progress[64] <= progress[63];
    always @(posedge clk) progress[65] <= progress[64];
    always @(posedge clk) progress[66] <= progress[65];
    always @(posedge clk) progress[67] <= progress[66];
    always @(posedge clk) progress[68] <= progress[67];
    always @(posedge clk) progress[69] <= progress[68];
    always @(posedge clk) progress[70] <= progress[69];
    always @(posedge clk) progress[71] <= progress[70];
    always @(posedge clk) progress[72] <= progress[71];
    always @(posedge clk) progress[73] <= progress[72];
    always @(posedge clk) progress[74] <= progress[73];
    always @(posedge clk) progress[75] <= progress[74];
    always @(posedge clk) progress[76] <= progress[75];
    always @(posedge clk) progress[77] <= progress[76];
    always @(posedge clk) progress[78] <= progress[77];
    always @(posedge clk) progress[79] <= progress[78];
    always @(posedge clk) progress[80] <= progress[79];
    always @(posedge clk) progress[81] <= progress[80];
    always @(posedge clk) progress[82] <= progress[81];
    always @(posedge clk) progress[83] <= progress[82];
    always @(posedge clk) progress[84] <= progress[83];
    always @(posedge clk) progress[85] <= progress[84];
    always @(posedge clk) progress[86] <= progress[85];
    always @(posedge clk) progress[87] <= progress[86];
    always @(posedge clk) progress[88] <= progress[87];
    always @(posedge clk) progress[89] <= progress[88];
    always @(posedge clk) progress[90] <= progress[89];
    always @(posedge clk) progress[91] <= progress[90];
    always @(posedge clk) progress[92] <= progress[91];
    always @(posedge clk) progress[93] <= progress[92];
    always @(posedge clk) progress[94] <= progress[93];
    always @(posedge clk) progress[95] <= progress[94];
    always @(posedge clk) progress[96] <= progress[95];
    always @(posedge clk) progress[97] <= progress[96];
    always @(posedge clk) progress[98] <= progress[97];
    always @(posedge clk) progress[99] <= progress[98];
    always @(posedge clk) progress[100] <= progress[99];
    always @(posedge clk) progress[101] <= progress[100];
    always @(posedge clk) progress[102] <= progress[101];
    always @(posedge clk) progress[103] <= progress[102];
    always @(posedge clk) progress[104] <= progress[103];
    always @(posedge clk) progress[105] <= progress[104];
    always @(posedge clk) progress[106] <= progress[105];
    always @(posedge clk) progress[107] <= progress[106];
    always @(posedge clk) progress[108] <= progress[107];
    always @(posedge clk) progress[109] <= progress[108];
    always @(posedge clk) progress[110] <= progress[109];
    always @(posedge clk) progress[111] <= progress[110];
    always @(posedge clk) progress[112] <= progress[111];
    always @(posedge clk) progress[113] <= progress[112];
    always @(posedge clk) progress[114] <= progress[113];
    always @(posedge clk) progress[115] <= progress[114];
    always @(posedge clk) progress[116] <= progress[115];
    always @(posedge clk) progress[117] <= progress[116];
    always @(posedge clk) progress[118] <= progress[117];
    always @(posedge clk) progress[119] <= progress[118];
    always @(posedge clk) progress[120] <= progress[119];
    always @(posedge clk) progress[121] <= progress[120];
    always @(posedge clk) progress[122] <= progress[121];
    always @(posedge clk) progress[123] <= progress[122];
    always @(posedge clk) progress[124] <= progress[123];
    always @(posedge clk) progress[125] <= progress[124];
    always @(posedge clk) progress[126] <= progress[125];
    always @(posedge clk) progress[127] <= progress[126];
    always @(posedge clk) progress[128] <= progress[127];
    always @(posedge clk) progress[129] <= progress[128];
    always @(posedge clk) progress[130] <= progress[129];
    always @(posedge clk) progress[131] <= progress[130];
    always @(posedge clk) progress[132] <= progress[131];
    always @(posedge clk) progress[133] <= progress[132];
    always @(posedge clk) progress[134] <= progress[133];
    always @(posedge clk) progress[135] <= progress[134];
    always @(posedge clk) progress[136] <= progress[135];
    always @(posedge clk) progress[137] <= progress[136];
    always @(posedge clk) progress[138] <= progress[137];
    always @(posedge clk) progress[139] <= progress[138];
    always @(posedge clk) progress[140] <= progress[139];
    always @(posedge clk) progress[141] <= progress[140];
    always @(posedge clk) progress[142] <= progress[141];
    always @(posedge clk) progress[143] <= progress[142];
    always @(posedge clk) progress[144] <= progress[143];
    always @(posedge clk) progress[145] <= progress[144];
    always @(posedge clk) progress[146] <= progress[145];
    always @(posedge clk) progress[147] <= progress[146];
    always @(posedge clk) progress[148] <= progress[147];
    always @(posedge clk) progress[149] <= progress[148];
    always @(posedge clk) progress[150] <= progress[149];
    always @(posedge clk) progress[151] <= progress[150];
    always @(posedge clk) progress[152] <= progress[151];
    always @(posedge clk) progress[153] <= progress[152];
    always @(posedge clk) progress[154] <= progress[153];
    always @(posedge clk) progress[155] <= progress[154];
    always @(posedge clk) progress[156] <= progress[155];
    always @(posedge clk) progress[157] <= progress[156];
    always @(posedge clk) progress[158] <= progress[157];
    always @(posedge clk) progress[159] <= progress[158];
    always @(posedge clk) progress[160] <= progress[159];
    always @(posedge clk) progress[161] <= progress[160];
    always @(posedge clk) progress[162] <= progress[161];
    always @(posedge clk) progress[163] <= progress[162];
    always @(posedge clk) progress[164] <= progress[163];
    always @(posedge clk) progress[165] <= progress[164];
    always @(posedge clk) progress[166] <= progress[165];
    always @(posedge clk) progress[167] <= progress[166];
    always @(posedge clk) progress[168] <= progress[167];
    always @(posedge clk) progress[169] <= progress[168];
    always @(posedge clk) progress[170] <= progress[169];
    always @(posedge clk) progress[171] <= progress[170];
    always @(posedge clk) progress[172] <= progress[171];
    always @(posedge clk) progress[173] <= progress[172];
    always @(posedge clk) progress[174] <= progress[173];
    always @(posedge clk) progress[175] <= progress[174];
    always @(posedge clk) progress[176] <= progress[175];
    always @(posedge clk) progress[177] <= progress[176];
    assign write = progress[177];
endmodule

