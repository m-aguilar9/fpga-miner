module odo_pre_mix(in, out);
    input [639:0] in;
    output [639:0] out;
    wire [63:0] total;
    assign total = 0 ^ in[63:0] ^ in[127:64] ^ in[191:128] ^ in[255:192] ^ in[319:256] ^ in[383:320] ^ in[447:384] ^ in[511:448] ^ in[575:512] ^ in[639:576];
    assign out[63:0] = in[63:0] ^ total ^ (total >> 32);
    assign out[127:64] = in[127:64] ^ total ^ (total >> 32);
    assign out[191:128] = in[191:128] ^ total ^ (total >> 32);
    assign out[255:192] = in[255:192] ^ total ^ (total >> 32);
    assign out[319:256] = in[319:256] ^ total ^ (total >> 32);
    assign out[383:320] = in[383:320] ^ total ^ (total >> 32);
    assign out[447:384] = in[447:384] ^ total ^ (total >> 32);
    assign out[511:448] = in[511:448] ^ total ^ (total >> 32);
    assign out[575:512] = in[575:512] ^ total ^ (total >> 32);
    assign out[639:576] = in[639:576] ^ total ^ (total >> 32);
endmodule

module odo_sbox_small0(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h28;
        mem[1] = 6'h10;
        mem[2] = 6'h34;
        mem[3] = 6'h31;
        mem[4] = 6'h01;
        mem[5] = 6'h03;
        mem[6] = 6'h04;
        mem[7] = 6'h24;
        mem[8] = 6'h1b;
        mem[9] = 6'h33;
        mem[10] = 6'h1a;
        mem[11] = 6'h0e;
        mem[12] = 6'h2d;
        mem[13] = 6'h3e;
        mem[14] = 6'h07;
        mem[15] = 6'h3a;
        mem[16] = 6'h1e;
        mem[17] = 6'h02;
        mem[18] = 6'h13;
        mem[19] = 6'h05;
        mem[20] = 6'h1c;
        mem[21] = 6'h17;
        mem[22] = 6'h18;
        mem[23] = 6'h3d;
        mem[24] = 6'h09;
        mem[25] = 6'h2b;
        mem[26] = 6'h2f;
        mem[27] = 6'h0b;
        mem[28] = 6'h37;
        mem[29] = 6'h3b;
        mem[30] = 6'h0f;
        mem[31] = 6'h3c;
        mem[32] = 6'h23;
        mem[33] = 6'h14;
        mem[34] = 6'h15;
        mem[35] = 6'h29;
        mem[36] = 6'h16;
        mem[37] = 6'h3f;
        mem[38] = 6'h0d;
        mem[39] = 6'h22;
        mem[40] = 6'h39;
        mem[41] = 6'h11;
        mem[42] = 6'h2a;
        mem[43] = 6'h27;
        mem[44] = 6'h06;
        mem[45] = 6'h1d;
        mem[46] = 6'h38;
        mem[47] = 6'h19;
        mem[48] = 6'h0a;
        mem[49] = 6'h1f;
        mem[50] = 6'h0c;
        mem[51] = 6'h12;
        mem[52] = 6'h08;
        mem[53] = 6'h35;
        mem[54] = 6'h00;
        mem[55] = 6'h21;
        mem[56] = 6'h25;
        mem[57] = 6'h2c;
        mem[58] = 6'h36;
        mem[59] = 6'h20;
        mem[60] = 6'h30;
        mem[61] = 6'h32;
        mem[62] = 6'h26;
        mem[63] = 6'h2e;
    end
endmodule

module odo_sbox_small1(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h34;
        mem[1] = 6'h37;
        mem[2] = 6'h23;
        mem[3] = 6'h10;
        mem[4] = 6'h03;
        mem[5] = 6'h06;
        mem[6] = 6'h12;
        mem[7] = 6'h3b;
        mem[8] = 6'h1f;
        mem[9] = 6'h11;
        mem[10] = 6'h1e;
        mem[11] = 6'h28;
        mem[12] = 6'h39;
        mem[13] = 6'h0b;
        mem[14] = 6'h2c;
        mem[15] = 6'h0f;
        mem[16] = 6'h26;
        mem[17] = 6'h05;
        mem[18] = 6'h0a;
        mem[19] = 6'h24;
        mem[20] = 6'h22;
        mem[21] = 6'h0d;
        mem[22] = 6'h1c;
        mem[23] = 6'h04;
        mem[24] = 6'h14;
        mem[25] = 6'h3f;
        mem[26] = 6'h00;
        mem[27] = 6'h3d;
        mem[28] = 6'h32;
        mem[29] = 6'h15;
        mem[30] = 6'h1d;
        mem[31] = 6'h33;
        mem[32] = 6'h2d;
        mem[33] = 6'h17;
        mem[34] = 6'h29;
        mem[35] = 6'h0c;
        mem[36] = 6'h02;
        mem[37] = 6'h09;
        mem[38] = 6'h31;
        mem[39] = 6'h20;
        mem[40] = 6'h36;
        mem[41] = 6'h3a;
        mem[42] = 6'h38;
        mem[43] = 6'h3c;
        mem[44] = 6'h0e;
        mem[45] = 6'h1b;
        mem[46] = 6'h13;
        mem[47] = 6'h1a;
        mem[48] = 6'h2a;
        mem[49] = 6'h07;
        mem[50] = 6'h2f;
        mem[51] = 6'h19;
        mem[52] = 6'h21;
        mem[53] = 6'h01;
        mem[54] = 6'h16;
        mem[55] = 6'h08;
        mem[56] = 6'h35;
        mem[57] = 6'h18;
        mem[58] = 6'h30;
        mem[59] = 6'h2e;
        mem[60] = 6'h25;
        mem[61] = 6'h27;
        mem[62] = 6'h3e;
        mem[63] = 6'h2b;
    end
endmodule

module odo_sbox_small2(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h20;
        mem[1] = 6'h2f;
        mem[2] = 6'h1c;
        mem[3] = 6'h37;
        mem[4] = 6'h03;
        mem[5] = 6'h0b;
        mem[6] = 6'h19;
        mem[7] = 6'h04;
        mem[8] = 6'h0d;
        mem[9] = 6'h3b;
        mem[10] = 6'h02;
        mem[11] = 6'h25;
        mem[12] = 6'h05;
        mem[13] = 6'h21;
        mem[14] = 6'h13;
        mem[15] = 6'h3a;
        mem[16] = 6'h3c;
        mem[17] = 6'h0a;
        mem[18] = 6'h12;
        mem[19] = 6'h1b;
        mem[20] = 6'h2a;
        mem[21] = 6'h28;
        mem[22] = 6'h1f;
        mem[23] = 6'h34;
        mem[24] = 6'h2c;
        mem[25] = 6'h2d;
        mem[26] = 6'h0f;
        mem[27] = 6'h24;
        mem[28] = 6'h38;
        mem[29] = 6'h3d;
        mem[30] = 6'h1d;
        mem[31] = 6'h22;
        mem[32] = 6'h31;
        mem[33] = 6'h0c;
        mem[34] = 6'h09;
        mem[35] = 6'h33;
        mem[36] = 6'h00;
        mem[37] = 6'h30;
        mem[38] = 6'h3f;
        mem[39] = 6'h29;
        mem[40] = 6'h36;
        mem[41] = 6'h26;
        mem[42] = 6'h35;
        mem[43] = 6'h2b;
        mem[44] = 6'h17;
        mem[45] = 6'h08;
        mem[46] = 6'h07;
        mem[47] = 6'h1a;
        mem[48] = 6'h39;
        mem[49] = 6'h10;
        mem[50] = 6'h18;
        mem[51] = 6'h01;
        mem[52] = 6'h32;
        mem[53] = 6'h11;
        mem[54] = 6'h27;
        mem[55] = 6'h1e;
        mem[56] = 6'h2e;
        mem[57] = 6'h15;
        mem[58] = 6'h23;
        mem[59] = 6'h16;
        mem[60] = 6'h0e;
        mem[61] = 6'h14;
        mem[62] = 6'h3e;
        mem[63] = 6'h06;
    end
endmodule

module odo_sbox_small3(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3b;
        mem[1] = 6'h3c;
        mem[2] = 6'h15;
        mem[3] = 6'h21;
        mem[4] = 6'h1f;
        mem[5] = 6'h2d;
        mem[6] = 6'h38;
        mem[7] = 6'h0a;
        mem[8] = 6'h23;
        mem[9] = 6'h25;
        mem[10] = 6'h18;
        mem[11] = 6'h37;
        mem[12] = 6'h17;
        mem[13] = 6'h36;
        mem[14] = 6'h3f;
        mem[15] = 6'h31;
        mem[16] = 6'h05;
        mem[17] = 6'h01;
        mem[18] = 6'h27;
        mem[19] = 6'h2a;
        mem[20] = 6'h04;
        mem[21] = 6'h2f;
        mem[22] = 6'h2e;
        mem[23] = 6'h07;
        mem[24] = 6'h33;
        mem[25] = 6'h08;
        mem[26] = 6'h39;
        mem[27] = 6'h11;
        mem[28] = 6'h3d;
        mem[29] = 6'h1e;
        mem[30] = 6'h34;
        mem[31] = 6'h3e;
        mem[32] = 6'h12;
        mem[33] = 6'h00;
        mem[34] = 6'h10;
        mem[35] = 6'h24;
        mem[36] = 6'h20;
        mem[37] = 6'h1b;
        mem[38] = 6'h0f;
        mem[39] = 6'h02;
        mem[40] = 6'h29;
        mem[41] = 6'h3a;
        mem[42] = 6'h0b;
        mem[43] = 6'h13;
        mem[44] = 6'h0c;
        mem[45] = 6'h19;
        mem[46] = 6'h1a;
        mem[47] = 6'h06;
        mem[48] = 6'h0d;
        mem[49] = 6'h14;
        mem[50] = 6'h26;
        mem[51] = 6'h2c;
        mem[52] = 6'h2b;
        mem[53] = 6'h1c;
        mem[54] = 6'h0e;
        mem[55] = 6'h32;
        mem[56] = 6'h03;
        mem[57] = 6'h35;
        mem[58] = 6'h22;
        mem[59] = 6'h09;
        mem[60] = 6'h1d;
        mem[61] = 6'h30;
        mem[62] = 6'h16;
        mem[63] = 6'h28;
    end
endmodule

module odo_sbox_small4(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1c;
        mem[1] = 6'h07;
        mem[2] = 6'h22;
        mem[3] = 6'h2a;
        mem[4] = 6'h29;
        mem[5] = 6'h32;
        mem[6] = 6'h02;
        mem[7] = 6'h03;
        mem[8] = 6'h2e;
        mem[9] = 6'h18;
        mem[10] = 6'h0b;
        mem[11] = 6'h0c;
        mem[12] = 6'h1b;
        mem[13] = 6'h26;
        mem[14] = 6'h0e;
        mem[15] = 6'h1d;
        mem[16] = 6'h16;
        mem[17] = 6'h28;
        mem[18] = 6'h27;
        mem[19] = 6'h30;
        mem[20] = 6'h38;
        mem[21] = 6'h12;
        mem[22] = 6'h33;
        mem[23] = 6'h25;
        mem[24] = 6'h17;
        mem[25] = 6'h13;
        mem[26] = 6'h21;
        mem[27] = 6'h1a;
        mem[28] = 6'h01;
        mem[29] = 6'h3d;
        mem[30] = 6'h24;
        mem[31] = 6'h05;
        mem[32] = 6'h10;
        mem[33] = 6'h08;
        mem[34] = 6'h2d;
        mem[35] = 6'h3f;
        mem[36] = 6'h3b;
        mem[37] = 6'h23;
        mem[38] = 6'h0d;
        mem[39] = 6'h11;
        mem[40] = 6'h1f;
        mem[41] = 6'h3e;
        mem[42] = 6'h04;
        mem[43] = 6'h00;
        mem[44] = 6'h09;
        mem[45] = 6'h0f;
        mem[46] = 6'h35;
        mem[47] = 6'h31;
        mem[48] = 6'h3a;
        mem[49] = 6'h2c;
        mem[50] = 6'h20;
        mem[51] = 6'h1e;
        mem[52] = 6'h19;
        mem[53] = 6'h36;
        mem[54] = 6'h37;
        mem[55] = 6'h0a;
        mem[56] = 6'h34;
        mem[57] = 6'h39;
        mem[58] = 6'h15;
        mem[59] = 6'h06;
        mem[60] = 6'h14;
        mem[61] = 6'h3c;
        mem[62] = 6'h2b;
        mem[63] = 6'h2f;
    end
endmodule

module odo_sbox_small5(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0e;
        mem[1] = 6'h13;
        mem[2] = 6'h3f;
        mem[3] = 6'h38;
        mem[4] = 6'h1c;
        mem[5] = 6'h08;
        mem[6] = 6'h3d;
        mem[7] = 6'h21;
        mem[8] = 6'h16;
        mem[9] = 6'h20;
        mem[10] = 6'h28;
        mem[11] = 6'h1a;
        mem[12] = 6'h33;
        mem[13] = 6'h11;
        mem[14] = 6'h22;
        mem[15] = 6'h17;
        mem[16] = 6'h00;
        mem[17] = 6'h1b;
        mem[18] = 6'h04;
        mem[19] = 6'h23;
        mem[20] = 6'h10;
        mem[21] = 6'h35;
        mem[22] = 6'h30;
        mem[23] = 6'h02;
        mem[24] = 6'h2d;
        mem[25] = 6'h24;
        mem[26] = 6'h01;
        mem[27] = 6'h03;
        mem[28] = 6'h18;
        mem[29] = 6'h3c;
        mem[30] = 6'h15;
        mem[31] = 6'h27;
        mem[32] = 6'h06;
        mem[33] = 6'h2f;
        mem[34] = 6'h1d;
        mem[35] = 6'h25;
        mem[36] = 6'h3a;
        mem[37] = 6'h0a;
        mem[38] = 6'h29;
        mem[39] = 6'h19;
        mem[40] = 6'h0b;
        mem[41] = 6'h32;
        mem[42] = 6'h05;
        mem[43] = 6'h36;
        mem[44] = 6'h3e;
        mem[45] = 6'h0c;
        mem[46] = 6'h0f;
        mem[47] = 6'h26;
        mem[48] = 6'h2a;
        mem[49] = 6'h1f;
        mem[50] = 6'h1e;
        mem[51] = 6'h14;
        mem[52] = 6'h3b;
        mem[53] = 6'h2e;
        mem[54] = 6'h0d;
        mem[55] = 6'h39;
        mem[56] = 6'h09;
        mem[57] = 6'h34;
        mem[58] = 6'h2b;
        mem[59] = 6'h12;
        mem[60] = 6'h2c;
        mem[61] = 6'h37;
        mem[62] = 6'h31;
        mem[63] = 6'h07;
    end
endmodule

module odo_sbox_small6(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1e;
        mem[1] = 6'h30;
        mem[2] = 6'h26;
        mem[3] = 6'h28;
        mem[4] = 6'h3d;
        mem[5] = 6'h37;
        mem[6] = 6'h19;
        mem[7] = 6'h3e;
        mem[8] = 6'h38;
        mem[9] = 6'h13;
        mem[10] = 6'h10;
        mem[11] = 6'h0c;
        mem[12] = 6'h1f;
        mem[13] = 6'h05;
        mem[14] = 6'h16;
        mem[15] = 6'h03;
        mem[16] = 6'h15;
        mem[17] = 6'h1a;
        mem[18] = 6'h01;
        mem[19] = 6'h0b;
        mem[20] = 6'h2a;
        mem[21] = 6'h1c;
        mem[22] = 6'h07;
        mem[23] = 6'h33;
        mem[24] = 6'h02;
        mem[25] = 6'h3b;
        mem[26] = 6'h20;
        mem[27] = 6'h34;
        mem[28] = 6'h06;
        mem[29] = 6'h00;
        mem[30] = 6'h2e;
        mem[31] = 6'h2d;
        mem[32] = 6'h3c;
        mem[33] = 6'h08;
        mem[34] = 6'h04;
        mem[35] = 6'h3a;
        mem[36] = 6'h17;
        mem[37] = 6'h23;
        mem[38] = 6'h27;
        mem[39] = 6'h1b;
        mem[40] = 6'h1d;
        mem[41] = 6'h12;
        mem[42] = 6'h29;
        mem[43] = 6'h35;
        mem[44] = 6'h0d;
        mem[45] = 6'h14;
        mem[46] = 6'h22;
        mem[47] = 6'h18;
        mem[48] = 6'h24;
        mem[49] = 6'h11;
        mem[50] = 6'h36;
        mem[51] = 6'h39;
        mem[52] = 6'h32;
        mem[53] = 6'h2f;
        mem[54] = 6'h21;
        mem[55] = 6'h3f;
        mem[56] = 6'h25;
        mem[57] = 6'h0a;
        mem[58] = 6'h0e;
        mem[59] = 6'h31;
        mem[60] = 6'h0f;
        mem[61] = 6'h09;
        mem[62] = 6'h2c;
        mem[63] = 6'h2b;
    end
endmodule

module odo_sbox_small7(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h19;
        mem[1] = 6'h0d;
        mem[2] = 6'h3e;
        mem[3] = 6'h36;
        mem[4] = 6'h0c;
        mem[5] = 6'h2c;
        mem[6] = 6'h13;
        mem[7] = 6'h3b;
        mem[8] = 6'h00;
        mem[9] = 6'h27;
        mem[10] = 6'h2e;
        mem[11] = 6'h0e;
        mem[12] = 6'h3f;
        mem[13] = 6'h07;
        mem[14] = 6'h3d;
        mem[15] = 6'h32;
        mem[16] = 6'h3a;
        mem[17] = 6'h22;
        mem[18] = 6'h35;
        mem[19] = 6'h24;
        mem[20] = 6'h26;
        mem[21] = 6'h3c;
        mem[22] = 6'h1a;
        mem[23] = 6'h28;
        mem[24] = 6'h25;
        mem[25] = 6'h0b;
        mem[26] = 6'h33;
        mem[27] = 6'h39;
        mem[28] = 6'h0f;
        mem[29] = 6'h29;
        mem[30] = 6'h20;
        mem[31] = 6'h34;
        mem[32] = 6'h21;
        mem[33] = 6'h08;
        mem[34] = 6'h23;
        mem[35] = 6'h2b;
        mem[36] = 6'h06;
        mem[37] = 6'h1c;
        mem[38] = 6'h1b;
        mem[39] = 6'h16;
        mem[40] = 6'h38;
        mem[41] = 6'h2d;
        mem[42] = 6'h11;
        mem[43] = 6'h18;
        mem[44] = 6'h2a;
        mem[45] = 6'h1e;
        mem[46] = 6'h04;
        mem[47] = 6'h2f;
        mem[48] = 6'h1f;
        mem[49] = 6'h30;
        mem[50] = 6'h09;
        mem[51] = 6'h10;
        mem[52] = 6'h01;
        mem[53] = 6'h14;
        mem[54] = 6'h37;
        mem[55] = 6'h1d;
        mem[56] = 6'h03;
        mem[57] = 6'h05;
        mem[58] = 6'h02;
        mem[59] = 6'h31;
        mem[60] = 6'h0a;
        mem[61] = 6'h15;
        mem[62] = 6'h17;
        mem[63] = 6'h12;
    end
endmodule

module odo_sbox_small8(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h05;
        mem[1] = 6'h2a;
        mem[2] = 6'h03;
        mem[3] = 6'h07;
        mem[4] = 6'h0f;
        mem[5] = 6'h3c;
        mem[6] = 6'h3e;
        mem[7] = 6'h08;
        mem[8] = 6'h33;
        mem[9] = 6'h0b;
        mem[10] = 6'h3d;
        mem[11] = 6'h14;
        mem[12] = 6'h0a;
        mem[13] = 6'h15;
        mem[14] = 6'h35;
        mem[15] = 6'h24;
        mem[16] = 6'h20;
        mem[17] = 6'h1b;
        mem[18] = 6'h13;
        mem[19] = 6'h38;
        mem[20] = 6'h1d;
        mem[21] = 6'h10;
        mem[22] = 6'h34;
        mem[23] = 6'h32;
        mem[24] = 6'h04;
        mem[25] = 6'h22;
        mem[26] = 6'h39;
        mem[27] = 6'h0d;
        mem[28] = 6'h2c;
        mem[29] = 6'h16;
        mem[30] = 6'h1e;
        mem[31] = 6'h3f;
        mem[32] = 6'h17;
        mem[33] = 6'h00;
        mem[34] = 6'h28;
        mem[35] = 6'h26;
        mem[36] = 6'h2e;
        mem[37] = 6'h06;
        mem[38] = 6'h12;
        mem[39] = 6'h0c;
        mem[40] = 6'h29;
        mem[41] = 6'h2d;
        mem[42] = 6'h1a;
        mem[43] = 6'h27;
        mem[44] = 6'h3a;
        mem[45] = 6'h3b;
        mem[46] = 6'h30;
        mem[47] = 6'h11;
        mem[48] = 6'h1f;
        mem[49] = 6'h37;
        mem[50] = 6'h36;
        mem[51] = 6'h01;
        mem[52] = 6'h25;
        mem[53] = 6'h2f;
        mem[54] = 6'h02;
        mem[55] = 6'h1c;
        mem[56] = 6'h23;
        mem[57] = 6'h19;
        mem[58] = 6'h18;
        mem[59] = 6'h31;
        mem[60] = 6'h21;
        mem[61] = 6'h09;
        mem[62] = 6'h2b;
        mem[63] = 6'h0e;
    end
endmodule

module odo_sbox_small9(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2d;
        mem[1] = 6'h19;
        mem[2] = 6'h25;
        mem[3] = 6'h33;
        mem[4] = 6'h1e;
        mem[5] = 6'h32;
        mem[6] = 6'h38;
        mem[7] = 6'h1c;
        mem[8] = 6'h22;
        mem[9] = 6'h06;
        mem[10] = 6'h2c;
        mem[11] = 6'h36;
        mem[12] = 6'h03;
        mem[13] = 6'h1b;
        mem[14] = 6'h07;
        mem[15] = 6'h1f;
        mem[16] = 6'h11;
        mem[17] = 6'h15;
        mem[18] = 6'h0d;
        mem[19] = 6'h28;
        mem[20] = 6'h17;
        mem[21] = 6'h3d;
        mem[22] = 6'h23;
        mem[23] = 6'h2e;
        mem[24] = 6'h3e;
        mem[25] = 6'h30;
        mem[26] = 6'h29;
        mem[27] = 6'h18;
        mem[28] = 6'h00;
        mem[29] = 6'h37;
        mem[30] = 6'h0a;
        mem[31] = 6'h0c;
        mem[32] = 6'h0f;
        mem[33] = 6'h0b;
        mem[34] = 6'h13;
        mem[35] = 6'h26;
        mem[36] = 6'h14;
        mem[37] = 6'h05;
        mem[38] = 6'h2a;
        mem[39] = 6'h01;
        mem[40] = 6'h0e;
        mem[41] = 6'h2b;
        mem[42] = 6'h31;
        mem[43] = 6'h02;
        mem[44] = 6'h3f;
        mem[45] = 6'h27;
        mem[46] = 6'h08;
        mem[47] = 6'h21;
        mem[48] = 6'h39;
        mem[49] = 6'h2f;
        mem[50] = 6'h16;
        mem[51] = 6'h3b;
        mem[52] = 6'h04;
        mem[53] = 6'h35;
        mem[54] = 6'h24;
        mem[55] = 6'h12;
        mem[56] = 6'h1d;
        mem[57] = 6'h20;
        mem[58] = 6'h3a;
        mem[59] = 6'h1a;
        mem[60] = 6'h3c;
        mem[61] = 6'h34;
        mem[62] = 6'h10;
        mem[63] = 6'h09;
    end
endmodule

module odo_sbox_small10(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2a;
        mem[1] = 6'h38;
        mem[2] = 6'h0e;
        mem[3] = 6'h2d;
        mem[4] = 6'h2e;
        mem[5] = 6'h2c;
        mem[6] = 6'h36;
        mem[7] = 6'h27;
        mem[8] = 6'h0a;
        mem[9] = 6'h1b;
        mem[10] = 6'h3e;
        mem[11] = 6'h14;
        mem[12] = 6'h3a;
        mem[13] = 6'h20;
        mem[14] = 6'h3b;
        mem[15] = 6'h3d;
        mem[16] = 6'h24;
        mem[17] = 6'h1d;
        mem[18] = 6'h09;
        mem[19] = 6'h05;
        mem[20] = 6'h2b;
        mem[21] = 6'h12;
        mem[22] = 6'h3c;
        mem[23] = 6'h0f;
        mem[24] = 6'h17;
        mem[25] = 6'h1f;
        mem[26] = 6'h10;
        mem[27] = 6'h3f;
        mem[28] = 6'h34;
        mem[29] = 6'h03;
        mem[30] = 6'h23;
        mem[31] = 6'h0d;
        mem[32] = 6'h04;
        mem[33] = 6'h26;
        mem[34] = 6'h08;
        mem[35] = 6'h11;
        mem[36] = 6'h0b;
        mem[37] = 6'h19;
        mem[38] = 6'h39;
        mem[39] = 6'h07;
        mem[40] = 6'h13;
        mem[41] = 6'h01;
        mem[42] = 6'h00;
        mem[43] = 6'h30;
        mem[44] = 6'h1a;
        mem[45] = 6'h25;
        mem[46] = 6'h21;
        mem[47] = 6'h02;
        mem[48] = 6'h33;
        mem[49] = 6'h28;
        mem[50] = 6'h31;
        mem[51] = 6'h0c;
        mem[52] = 6'h32;
        mem[53] = 6'h06;
        mem[54] = 6'h18;
        mem[55] = 6'h15;
        mem[56] = 6'h2f;
        mem[57] = 6'h37;
        mem[58] = 6'h22;
        mem[59] = 6'h35;
        mem[60] = 6'h1c;
        mem[61] = 6'h16;
        mem[62] = 6'h29;
        mem[63] = 6'h1e;
    end
endmodule

module odo_sbox_small11(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h03;
        mem[1] = 6'h23;
        mem[2] = 6'h29;
        mem[3] = 6'h35;
        mem[4] = 6'h1e;
        mem[5] = 6'h09;
        mem[6] = 6'h2b;
        mem[7] = 6'h3c;
        mem[8] = 6'h2e;
        mem[9] = 6'h19;
        mem[10] = 6'h25;
        mem[11] = 6'h2d;
        mem[12] = 6'h13;
        mem[13] = 6'h34;
        mem[14] = 6'h07;
        mem[15] = 6'h31;
        mem[16] = 6'h30;
        mem[17] = 6'h04;
        mem[18] = 6'h0b;
        mem[19] = 6'h21;
        mem[20] = 6'h06;
        mem[21] = 6'h37;
        mem[22] = 6'h1a;
        mem[23] = 6'h22;
        mem[24] = 6'h24;
        mem[25] = 6'h1c;
        mem[26] = 6'h16;
        mem[27] = 6'h00;
        mem[28] = 6'h01;
        mem[29] = 6'h10;
        mem[30] = 6'h08;
        mem[31] = 6'h15;
        mem[32] = 6'h3e;
        mem[33] = 6'h18;
        mem[34] = 6'h0a;
        mem[35] = 6'h0e;
        mem[36] = 6'h0d;
        mem[37] = 6'h3a;
        mem[38] = 6'h14;
        mem[39] = 6'h1f;
        mem[40] = 6'h0f;
        mem[41] = 6'h39;
        mem[42] = 6'h33;
        mem[43] = 6'h1b;
        mem[44] = 6'h11;
        mem[45] = 6'h12;
        mem[46] = 6'h02;
        mem[47] = 6'h3f;
        mem[48] = 6'h27;
        mem[49] = 6'h28;
        mem[50] = 6'h26;
        mem[51] = 6'h36;
        mem[52] = 6'h2a;
        mem[53] = 6'h2f;
        mem[54] = 6'h05;
        mem[55] = 6'h32;
        mem[56] = 6'h3b;
        mem[57] = 6'h20;
        mem[58] = 6'h1d;
        mem[59] = 6'h3d;
        mem[60] = 6'h38;
        mem[61] = 6'h2c;
        mem[62] = 6'h17;
        mem[63] = 6'h0c;
    end
endmodule

module odo_sbox_small12(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h23;
        mem[1] = 6'h24;
        mem[2] = 6'h17;
        mem[3] = 6'h06;
        mem[4] = 6'h25;
        mem[5] = 6'h1b;
        mem[6] = 6'h15;
        mem[7] = 6'h3b;
        mem[8] = 6'h0d;
        mem[9] = 6'h07;
        mem[10] = 6'h1e;
        mem[11] = 6'h1d;
        mem[12] = 6'h00;
        mem[13] = 6'h04;
        mem[14] = 6'h28;
        mem[15] = 6'h21;
        mem[16] = 6'h11;
        mem[17] = 6'h2d;
        mem[18] = 6'h0b;
        mem[19] = 6'h09;
        mem[20] = 6'h01;
        mem[21] = 6'h2a;
        mem[22] = 6'h34;
        mem[23] = 6'h0f;
        mem[24] = 6'h08;
        mem[25] = 6'h22;
        mem[26] = 6'h1f;
        mem[27] = 6'h2e;
        mem[28] = 6'h33;
        mem[29] = 6'h3e;
        mem[30] = 6'h35;
        mem[31] = 6'h13;
        mem[32] = 6'h1a;
        mem[33] = 6'h30;
        mem[34] = 6'h16;
        mem[35] = 6'h27;
        mem[36] = 6'h14;
        mem[37] = 6'h19;
        mem[38] = 6'h2f;
        mem[39] = 6'h36;
        mem[40] = 6'h20;
        mem[41] = 6'h02;
        mem[42] = 6'h3a;
        mem[43] = 6'h0c;
        mem[44] = 6'h03;
        mem[45] = 6'h32;
        mem[46] = 6'h2c;
        mem[47] = 6'h18;
        mem[48] = 6'h3c;
        mem[49] = 6'h37;
        mem[50] = 6'h05;
        mem[51] = 6'h26;
        mem[52] = 6'h29;
        mem[53] = 6'h2b;
        mem[54] = 6'h3d;
        mem[55] = 6'h1c;
        mem[56] = 6'h31;
        mem[57] = 6'h0e;
        mem[58] = 6'h0a;
        mem[59] = 6'h39;
        mem[60] = 6'h12;
        mem[61] = 6'h10;
        mem[62] = 6'h38;
        mem[63] = 6'h3f;
    end
endmodule

module odo_sbox_small13(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h04;
        mem[1] = 6'h01;
        mem[2] = 6'h3c;
        mem[3] = 6'h2c;
        mem[4] = 6'h1d;
        mem[5] = 6'h2b;
        mem[6] = 6'h09;
        mem[7] = 6'h19;
        mem[8] = 6'h1a;
        mem[9] = 6'h20;
        mem[10] = 6'h13;
        mem[11] = 6'h3d;
        mem[12] = 6'h3e;
        mem[13] = 6'h15;
        mem[14] = 6'h24;
        mem[15] = 6'h36;
        mem[16] = 6'h23;
        mem[17] = 6'h3f;
        mem[18] = 6'h2a;
        mem[19] = 6'h33;
        mem[20] = 6'h26;
        mem[21] = 6'h35;
        mem[22] = 6'h16;
        mem[23] = 6'h07;
        mem[24] = 6'h2f;
        mem[25] = 6'h1c;
        mem[26] = 6'h2e;
        mem[27] = 6'h22;
        mem[28] = 6'h1f;
        mem[29] = 6'h02;
        mem[30] = 6'h32;
        mem[31] = 6'h08;
        mem[32] = 6'h0a;
        mem[33] = 6'h1e;
        mem[34] = 6'h05;
        mem[35] = 6'h0d;
        mem[36] = 6'h00;
        mem[37] = 6'h3a;
        mem[38] = 6'h28;
        mem[39] = 6'h3b;
        mem[40] = 6'h18;
        mem[41] = 6'h38;
        mem[42] = 6'h0b;
        mem[43] = 6'h29;
        mem[44] = 6'h27;
        mem[45] = 6'h30;
        mem[46] = 6'h0f;
        mem[47] = 6'h37;
        mem[48] = 6'h03;
        mem[49] = 6'h0c;
        mem[50] = 6'h21;
        mem[51] = 6'h1b;
        mem[52] = 6'h06;
        mem[53] = 6'h39;
        mem[54] = 6'h14;
        mem[55] = 6'h25;
        mem[56] = 6'h11;
        mem[57] = 6'h34;
        mem[58] = 6'h10;
        mem[59] = 6'h12;
        mem[60] = 6'h0e;
        mem[61] = 6'h2d;
        mem[62] = 6'h17;
        mem[63] = 6'h31;
    end
endmodule

module odo_sbox_small14(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2b;
        mem[1] = 6'h39;
        mem[2] = 6'h1d;
        mem[3] = 6'h0f;
        mem[4] = 6'h2c;
        mem[5] = 6'h3b;
        mem[6] = 6'h3a;
        mem[7] = 6'h14;
        mem[8] = 6'h35;
        mem[9] = 6'h0a;
        mem[10] = 6'h37;
        mem[11] = 6'h30;
        mem[12] = 6'h09;
        mem[13] = 6'h11;
        mem[14] = 6'h25;
        mem[15] = 6'h21;
        mem[16] = 6'h23;
        mem[17] = 6'h17;
        mem[18] = 6'h22;
        mem[19] = 6'h1b;
        mem[20] = 6'h01;
        mem[21] = 6'h19;
        mem[22] = 6'h2a;
        mem[23] = 6'h00;
        mem[24] = 6'h05;
        mem[25] = 6'h2d;
        mem[26] = 6'h0c;
        mem[27] = 6'h1c;
        mem[28] = 6'h32;
        mem[29] = 6'h06;
        mem[30] = 6'h2f;
        mem[31] = 6'h38;
        mem[32] = 6'h33;
        mem[33] = 6'h34;
        mem[34] = 6'h02;
        mem[35] = 6'h1f;
        mem[36] = 6'h0d;
        mem[37] = 6'h18;
        mem[38] = 6'h16;
        mem[39] = 6'h15;
        mem[40] = 6'h3f;
        mem[41] = 6'h31;
        mem[42] = 6'h0b;
        mem[43] = 6'h10;
        mem[44] = 6'h3c;
        mem[45] = 6'h3d;
        mem[46] = 6'h04;
        mem[47] = 6'h3e;
        mem[48] = 6'h36;
        mem[49] = 6'h1a;
        mem[50] = 6'h29;
        mem[51] = 6'h0e;
        mem[52] = 6'h2e;
        mem[53] = 6'h03;
        mem[54] = 6'h28;
        mem[55] = 6'h20;
        mem[56] = 6'h26;
        mem[57] = 6'h07;
        mem[58] = 6'h1e;
        mem[59] = 6'h12;
        mem[60] = 6'h27;
        mem[61] = 6'h13;
        mem[62] = 6'h24;
        mem[63] = 6'h08;
    end
endmodule

module odo_sbox_small15(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2c;
        mem[1] = 6'h05;
        mem[2] = 6'h3e;
        mem[3] = 6'h34;
        mem[4] = 6'h0d;
        mem[5] = 6'h1a;
        mem[6] = 6'h28;
        mem[7] = 6'h38;
        mem[8] = 6'h20;
        mem[9] = 6'h12;
        mem[10] = 6'h0b;
        mem[11] = 6'h0c;
        mem[12] = 6'h2f;
        mem[13] = 6'h07;
        mem[14] = 6'h35;
        mem[15] = 6'h36;
        mem[16] = 6'h26;
        mem[17] = 6'h23;
        mem[18] = 6'h1e;
        mem[19] = 6'h1f;
        mem[20] = 6'h04;
        mem[21] = 6'h06;
        mem[22] = 6'h25;
        mem[23] = 6'h1b;
        mem[24] = 6'h2a;
        mem[25] = 6'h01;
        mem[26] = 6'h0a;
        mem[27] = 6'h17;
        mem[28] = 6'h30;
        mem[29] = 6'h31;
        mem[30] = 6'h3d;
        mem[31] = 6'h22;
        mem[32] = 6'h09;
        mem[33] = 6'h2d;
        mem[34] = 6'h16;
        mem[35] = 6'h19;
        mem[36] = 6'h18;
        mem[37] = 6'h2b;
        mem[38] = 6'h32;
        mem[39] = 6'h3b;
        mem[40] = 6'h3c;
        mem[41] = 6'h00;
        mem[42] = 6'h02;
        mem[43] = 6'h2e;
        mem[44] = 6'h29;
        mem[45] = 6'h21;
        mem[46] = 6'h37;
        mem[47] = 6'h10;
        mem[48] = 6'h3f;
        mem[49] = 6'h33;
        mem[50] = 6'h1d;
        mem[51] = 6'h1c;
        mem[52] = 6'h08;
        mem[53] = 6'h0e;
        mem[54] = 6'h24;
        mem[55] = 6'h14;
        mem[56] = 6'h0f;
        mem[57] = 6'h39;
        mem[58] = 6'h13;
        mem[59] = 6'h03;
        mem[60] = 6'h27;
        mem[61] = 6'h11;
        mem[62] = 6'h3a;
        mem[63] = 6'h15;
    end
endmodule

module odo_sbox_small16(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2c;
        mem[1] = 6'h38;
        mem[2] = 6'h30;
        mem[3] = 6'h3d;
        mem[4] = 6'h02;
        mem[5] = 6'h27;
        mem[6] = 6'h0e;
        mem[7] = 6'h22;
        mem[8] = 6'h0b;
        mem[9] = 6'h3b;
        mem[10] = 6'h17;
        mem[11] = 6'h25;
        mem[12] = 6'h16;
        mem[13] = 6'h2e;
        mem[14] = 6'h06;
        mem[15] = 6'h04;
        mem[16] = 6'h1a;
        mem[17] = 6'h09;
        mem[18] = 6'h32;
        mem[19] = 6'h19;
        mem[20] = 6'h1f;
        mem[21] = 6'h3f;
        mem[22] = 6'h21;
        mem[23] = 6'h2d;
        mem[24] = 6'h3e;
        mem[25] = 6'h1d;
        mem[26] = 6'h2a;
        mem[27] = 6'h3a;
        mem[28] = 6'h1c;
        mem[29] = 6'h0c;
        mem[30] = 6'h24;
        mem[31] = 6'h0a;
        mem[32] = 6'h11;
        mem[33] = 6'h0f;
        mem[34] = 6'h35;
        mem[35] = 6'h18;
        mem[36] = 6'h36;
        mem[37] = 6'h26;
        mem[38] = 6'h33;
        mem[39] = 6'h1e;
        mem[40] = 6'h37;
        mem[41] = 6'h1b;
        mem[42] = 6'h2b;
        mem[43] = 6'h0d;
        mem[44] = 6'h00;
        mem[45] = 6'h13;
        mem[46] = 6'h12;
        mem[47] = 6'h10;
        mem[48] = 6'h3c;
        mem[49] = 6'h2f;
        mem[50] = 6'h20;
        mem[51] = 6'h14;
        mem[52] = 6'h34;
        mem[53] = 6'h08;
        mem[54] = 6'h15;
        mem[55] = 6'h31;
        mem[56] = 6'h28;
        mem[57] = 6'h29;
        mem[58] = 6'h05;
        mem[59] = 6'h01;
        mem[60] = 6'h23;
        mem[61] = 6'h39;
        mem[62] = 6'h03;
        mem[63] = 6'h07;
    end
endmodule

module odo_sbox_small17(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h25;
        mem[1] = 6'h39;
        mem[2] = 6'h3c;
        mem[3] = 6'h3e;
        mem[4] = 6'h0c;
        mem[5] = 6'h21;
        mem[6] = 6'h27;
        mem[7] = 6'h20;
        mem[8] = 6'h14;
        mem[9] = 6'h08;
        mem[10] = 6'h13;
        mem[11] = 6'h2b;
        mem[12] = 6'h29;
        mem[13] = 6'h30;
        mem[14] = 6'h3f;
        mem[15] = 6'h2c;
        mem[16] = 6'h3b;
        mem[17] = 6'h38;
        mem[18] = 6'h3a;
        mem[19] = 6'h1d;
        mem[20] = 6'h37;
        mem[21] = 6'h26;
        mem[22] = 6'h12;
        mem[23] = 6'h02;
        mem[24] = 6'h05;
        mem[25] = 6'h1f;
        mem[26] = 6'h0f;
        mem[27] = 6'h31;
        mem[28] = 6'h22;
        mem[29] = 6'h15;
        mem[30] = 6'h16;
        mem[31] = 6'h0d;
        mem[32] = 6'h1a;
        mem[33] = 6'h19;
        mem[34] = 6'h3d;
        mem[35] = 6'h2d;
        mem[36] = 6'h01;
        mem[37] = 6'h34;
        mem[38] = 6'h0b;
        mem[39] = 6'h28;
        mem[40] = 6'h1c;
        mem[41] = 6'h36;
        mem[42] = 6'h0e;
        mem[43] = 6'h00;
        mem[44] = 6'h35;
        mem[45] = 6'h03;
        mem[46] = 6'h33;
        mem[47] = 6'h1b;
        mem[48] = 6'h07;
        mem[49] = 6'h04;
        mem[50] = 6'h24;
        mem[51] = 6'h2e;
        mem[52] = 6'h18;
        mem[53] = 6'h2a;
        mem[54] = 6'h06;
        mem[55] = 6'h2f;
        mem[56] = 6'h09;
        mem[57] = 6'h10;
        mem[58] = 6'h23;
        mem[59] = 6'h32;
        mem[60] = 6'h1e;
        mem[61] = 6'h0a;
        mem[62] = 6'h17;
        mem[63] = 6'h11;
    end
endmodule

module odo_sbox_small18(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h00;
        mem[1] = 6'h36;
        mem[2] = 6'h3d;
        mem[3] = 6'h0e;
        mem[4] = 6'h1d;
        mem[5] = 6'h05;
        mem[6] = 6'h12;
        mem[7] = 6'h07;
        mem[8] = 6'h1b;
        mem[9] = 6'h39;
        mem[10] = 6'h24;
        mem[11] = 6'h14;
        mem[12] = 6'h3c;
        mem[13] = 6'h2f;
        mem[14] = 6'h0f;
        mem[15] = 6'h17;
        mem[16] = 6'h18;
        mem[17] = 6'h0d;
        mem[18] = 6'h06;
        mem[19] = 6'h31;
        mem[20] = 6'h3a;
        mem[21] = 6'h25;
        mem[22] = 6'h2b;
        mem[23] = 6'h37;
        mem[24] = 6'h2a;
        mem[25] = 6'h1e;
        mem[26] = 6'h10;
        mem[27] = 6'h20;
        mem[28] = 6'h30;
        mem[29] = 6'h01;
        mem[30] = 6'h33;
        mem[31] = 6'h15;
        mem[32] = 6'h1c;
        mem[33] = 6'h23;
        mem[34] = 6'h35;
        mem[35] = 6'h34;
        mem[36] = 6'h11;
        mem[37] = 6'h22;
        mem[38] = 6'h02;
        mem[39] = 6'h08;
        mem[40] = 6'h13;
        mem[41] = 6'h1a;
        mem[42] = 6'h2c;
        mem[43] = 6'h38;
        mem[44] = 6'h26;
        mem[45] = 6'h2d;
        mem[46] = 6'h16;
        mem[47] = 6'h09;
        mem[48] = 6'h32;
        mem[49] = 6'h3f;
        mem[50] = 6'h0c;
        mem[51] = 6'h1f;
        mem[52] = 6'h27;
        mem[53] = 6'h3b;
        mem[54] = 6'h3e;
        mem[55] = 6'h21;
        mem[56] = 6'h2e;
        mem[57] = 6'h28;
        mem[58] = 6'h04;
        mem[59] = 6'h0a;
        mem[60] = 6'h0b;
        mem[61] = 6'h19;
        mem[62] = 6'h03;
        mem[63] = 6'h29;
    end
endmodule

module odo_sbox_small19(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h35;
        mem[1] = 6'h17;
        mem[2] = 6'h23;
        mem[3] = 6'h21;
        mem[4] = 6'h02;
        mem[5] = 6'h3f;
        mem[6] = 6'h19;
        mem[7] = 6'h18;
        mem[8] = 6'h00;
        mem[9] = 6'h12;
        mem[10] = 6'h30;
        mem[11] = 6'h36;
        mem[12] = 6'h15;
        mem[13] = 6'h33;
        mem[14] = 6'h06;
        mem[15] = 6'h1d;
        mem[16] = 6'h3e;
        mem[17] = 6'h2b;
        mem[18] = 6'h37;
        mem[19] = 6'h01;
        mem[20] = 6'h3c;
        mem[21] = 6'h04;
        mem[22] = 6'h0b;
        mem[23] = 6'h2e;
        mem[24] = 6'h3b;
        mem[25] = 6'h2d;
        mem[26] = 6'h2f;
        mem[27] = 6'h0c;
        mem[28] = 6'h1f;
        mem[29] = 6'h22;
        mem[30] = 6'h34;
        mem[31] = 6'h26;
        mem[32] = 6'h03;
        mem[33] = 6'h05;
        mem[34] = 6'h07;
        mem[35] = 6'h1a;
        mem[36] = 6'h0a;
        mem[37] = 6'h0e;
        mem[38] = 6'h14;
        mem[39] = 6'h25;
        mem[40] = 6'h1e;
        mem[41] = 6'h2a;
        mem[42] = 6'h3a;
        mem[43] = 6'h31;
        mem[44] = 6'h1c;
        mem[45] = 6'h09;
        mem[46] = 6'h13;
        mem[47] = 6'h39;
        mem[48] = 6'h32;
        mem[49] = 6'h2c;
        mem[50] = 6'h29;
        mem[51] = 6'h28;
        mem[52] = 6'h20;
        mem[53] = 6'h1b;
        mem[54] = 6'h24;
        mem[55] = 6'h38;
        mem[56] = 6'h16;
        mem[57] = 6'h0d;
        mem[58] = 6'h27;
        mem[59] = 6'h08;
        mem[60] = 6'h0f;
        mem[61] = 6'h10;
        mem[62] = 6'h3d;
        mem[63] = 6'h11;
    end
endmodule

module odo_sbox_small20(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h32;
        mem[1] = 6'h00;
        mem[2] = 6'h13;
        mem[3] = 6'h26;
        mem[4] = 6'h1d;
        mem[5] = 6'h28;
        mem[6] = 6'h2d;
        mem[7] = 6'h1c;
        mem[8] = 6'h38;
        mem[9] = 6'h18;
        mem[10] = 6'h3d;
        mem[11] = 6'h3c;
        mem[12] = 6'h05;
        mem[13] = 6'h1f;
        mem[14] = 6'h21;
        mem[15] = 6'h14;
        mem[16] = 6'h36;
        mem[17] = 6'h0e;
        mem[18] = 6'h25;
        mem[19] = 6'h3e;
        mem[20] = 6'h29;
        mem[21] = 6'h2c;
        mem[22] = 6'h35;
        mem[23] = 6'h0b;
        mem[24] = 6'h07;
        mem[25] = 6'h12;
        mem[26] = 6'h17;
        mem[27] = 6'h08;
        mem[28] = 6'h0d;
        mem[29] = 6'h30;
        mem[30] = 6'h37;
        mem[31] = 6'h33;
        mem[32] = 6'h10;
        mem[33] = 6'h39;
        mem[34] = 6'h01;
        mem[35] = 6'h22;
        mem[36] = 6'h24;
        mem[37] = 6'h1e;
        mem[38] = 6'h20;
        mem[39] = 6'h03;
        mem[40] = 6'h3a;
        mem[41] = 6'h2a;
        mem[42] = 6'h1a;
        mem[43] = 6'h3f;
        mem[44] = 6'h19;
        mem[45] = 6'h04;
        mem[46] = 6'h34;
        mem[47] = 6'h1b;
        mem[48] = 6'h23;
        mem[49] = 6'h2f;
        mem[50] = 6'h27;
        mem[51] = 6'h2e;
        mem[52] = 6'h02;
        mem[53] = 6'h06;
        mem[54] = 6'h09;
        mem[55] = 6'h16;
        mem[56] = 6'h31;
        mem[57] = 6'h0f;
        mem[58] = 6'h15;
        mem[59] = 6'h11;
        mem[60] = 6'h0c;
        mem[61] = 6'h3b;
        mem[62] = 6'h0a;
        mem[63] = 6'h2b;
    end
endmodule

module odo_sbox_small21(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h36;
        mem[1] = 6'h04;
        mem[2] = 6'h1d;
        mem[3] = 6'h2d;
        mem[4] = 6'h1b;
        mem[5] = 6'h2f;
        mem[6] = 6'h08;
        mem[7] = 6'h2e;
        mem[8] = 6'h3a;
        mem[9] = 6'h19;
        mem[10] = 6'h37;
        mem[11] = 6'h26;
        mem[12] = 6'h22;
        mem[13] = 6'h30;
        mem[14] = 6'h1f;
        mem[15] = 6'h29;
        mem[16] = 6'h38;
        mem[17] = 6'h24;
        mem[18] = 6'h23;
        mem[19] = 6'h06;
        mem[20] = 6'h13;
        mem[21] = 6'h0e;
        mem[22] = 6'h17;
        mem[23] = 6'h20;
        mem[24] = 6'h14;
        mem[25] = 6'h3f;
        mem[26] = 6'h12;
        mem[27] = 6'h32;
        mem[28] = 6'h16;
        mem[29] = 6'h09;
        mem[30] = 6'h0b;
        mem[31] = 6'h02;
        mem[32] = 6'h1a;
        mem[33] = 6'h34;
        mem[34] = 6'h2a;
        mem[35] = 6'h0f;
        mem[36] = 6'h00;
        mem[37] = 6'h15;
        mem[38] = 6'h25;
        mem[39] = 6'h39;
        mem[40] = 6'h03;
        mem[41] = 6'h3d;
        mem[42] = 6'h01;
        mem[43] = 6'h21;
        mem[44] = 6'h0d;
        mem[45] = 6'h3c;
        mem[46] = 6'h27;
        mem[47] = 6'h28;
        mem[48] = 6'h07;
        mem[49] = 6'h1c;
        mem[50] = 6'h0c;
        mem[51] = 6'h2c;
        mem[52] = 6'h10;
        mem[53] = 6'h0a;
        mem[54] = 6'h3b;
        mem[55] = 6'h11;
        mem[56] = 6'h31;
        mem[57] = 6'h05;
        mem[58] = 6'h18;
        mem[59] = 6'h33;
        mem[60] = 6'h3e;
        mem[61] = 6'h35;
        mem[62] = 6'h1e;
        mem[63] = 6'h2b;
    end
endmodule

module odo_sbox_small22(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h19;
        mem[1] = 6'h17;
        mem[2] = 6'h12;
        mem[3] = 6'h10;
        mem[4] = 6'h14;
        mem[5] = 6'h31;
        mem[6] = 6'h2c;
        mem[7] = 6'h2d;
        mem[8] = 6'h26;
        mem[9] = 6'h04;
        mem[10] = 6'h27;
        mem[11] = 6'h0a;
        mem[12] = 6'h3e;
        mem[13] = 6'h25;
        mem[14] = 6'h20;
        mem[15] = 6'h16;
        mem[16] = 6'h3a;
        mem[17] = 6'h09;
        mem[18] = 6'h0b;
        mem[19] = 6'h13;
        mem[20] = 6'h1f;
        mem[21] = 6'h1d;
        mem[22] = 6'h38;
        mem[23] = 6'h21;
        mem[24] = 6'h23;
        mem[25] = 6'h29;
        mem[26] = 6'h36;
        mem[27] = 6'h2b;
        mem[28] = 6'h07;
        mem[29] = 6'h0c;
        mem[30] = 6'h1c;
        mem[31] = 6'h1e;
        mem[32] = 6'h32;
        mem[33] = 6'h3b;
        mem[34] = 6'h08;
        mem[35] = 6'h2a;
        mem[36] = 6'h11;
        mem[37] = 6'h0f;
        mem[38] = 6'h2e;
        mem[39] = 6'h37;
        mem[40] = 6'h15;
        mem[41] = 6'h24;
        mem[42] = 6'h30;
        mem[43] = 6'h01;
        mem[44] = 6'h0e;
        mem[45] = 6'h28;
        mem[46] = 6'h22;
        mem[47] = 6'h06;
        mem[48] = 6'h2f;
        mem[49] = 6'h00;
        mem[50] = 6'h02;
        mem[51] = 6'h3f;
        mem[52] = 6'h33;
        mem[53] = 6'h0d;
        mem[54] = 6'h1a;
        mem[55] = 6'h3c;
        mem[56] = 6'h1b;
        mem[57] = 6'h34;
        mem[58] = 6'h3d;
        mem[59] = 6'h39;
        mem[60] = 6'h35;
        mem[61] = 6'h18;
        mem[62] = 6'h05;
        mem[63] = 6'h03;
    end
endmodule

module odo_sbox_small23(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0c;
        mem[1] = 6'h06;
        mem[2] = 6'h2f;
        mem[3] = 6'h34;
        mem[4] = 6'h36;
        mem[5] = 6'h38;
        mem[6] = 6'h3f;
        mem[7] = 6'h07;
        mem[8] = 6'h2c;
        mem[9] = 6'h27;
        mem[10] = 6'h16;
        mem[11] = 6'h3a;
        mem[12] = 6'h24;
        mem[13] = 6'h32;
        mem[14] = 6'h13;
        mem[15] = 6'h00;
        mem[16] = 6'h3c;
        mem[17] = 6'h31;
        mem[18] = 6'h02;
        mem[19] = 6'h12;
        mem[20] = 6'h15;
        mem[21] = 6'h20;
        mem[22] = 6'h2b;
        mem[23] = 6'h2a;
        mem[24] = 6'h1c;
        mem[25] = 6'h3d;
        mem[26] = 6'h03;
        mem[27] = 6'h23;
        mem[28] = 6'h1f;
        mem[29] = 6'h3b;
        mem[30] = 6'h10;
        mem[31] = 6'h21;
        mem[32] = 6'h1b;
        mem[33] = 6'h2e;
        mem[34] = 6'h39;
        mem[35] = 6'h01;
        mem[36] = 6'h37;
        mem[37] = 6'h18;
        mem[38] = 6'h17;
        mem[39] = 6'h14;
        mem[40] = 6'h0d;
        mem[41] = 6'h33;
        mem[42] = 6'h1a;
        mem[43] = 6'h1e;
        mem[44] = 6'h04;
        mem[45] = 6'h19;
        mem[46] = 6'h05;
        mem[47] = 6'h2d;
        mem[48] = 6'h28;
        mem[49] = 6'h22;
        mem[50] = 6'h0e;
        mem[51] = 6'h09;
        mem[52] = 6'h3e;
        mem[53] = 6'h0b;
        mem[54] = 6'h30;
        mem[55] = 6'h26;
        mem[56] = 6'h0a;
        mem[57] = 6'h1d;
        mem[58] = 6'h11;
        mem[59] = 6'h29;
        mem[60] = 6'h25;
        mem[61] = 6'h08;
        mem[62] = 6'h0f;
        mem[63] = 6'h35;
    end
endmodule

module odo_sbox_small24(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3a;
        mem[1] = 6'h06;
        mem[2] = 6'h0d;
        mem[3] = 6'h03;
        mem[4] = 6'h37;
        mem[5] = 6'h00;
        mem[6] = 6'h21;
        mem[7] = 6'h2c;
        mem[8] = 6'h38;
        mem[9] = 6'h11;
        mem[10] = 6'h26;
        mem[11] = 6'h08;
        mem[12] = 6'h2a;
        mem[13] = 6'h10;
        mem[14] = 6'h34;
        mem[15] = 6'h0f;
        mem[16] = 6'h16;
        mem[17] = 6'h3b;
        mem[18] = 6'h0a;
        mem[19] = 6'h02;
        mem[20] = 6'h19;
        mem[21] = 6'h3e;
        mem[22] = 6'h2f;
        mem[23] = 6'h0b;
        mem[24] = 6'h23;
        mem[25] = 6'h22;
        mem[26] = 6'h0e;
        mem[27] = 6'h2d;
        mem[28] = 6'h14;
        mem[29] = 6'h3c;
        mem[30] = 6'h32;
        mem[31] = 6'h3d;
        mem[32] = 6'h1b;
        mem[33] = 6'h29;
        mem[34] = 6'h25;
        mem[35] = 6'h13;
        mem[36] = 6'h18;
        mem[37] = 6'h36;
        mem[38] = 6'h33;
        mem[39] = 6'h05;
        mem[40] = 6'h1d;
        mem[41] = 6'h1e;
        mem[42] = 6'h24;
        mem[43] = 6'h04;
        mem[44] = 6'h30;
        mem[45] = 6'h35;
        mem[46] = 6'h01;
        mem[47] = 6'h3f;
        mem[48] = 6'h07;
        mem[49] = 6'h15;
        mem[50] = 6'h31;
        mem[51] = 6'h09;
        mem[52] = 6'h28;
        mem[53] = 6'h27;
        mem[54] = 6'h2e;
        mem[55] = 6'h0c;
        mem[56] = 6'h12;
        mem[57] = 6'h1a;
        mem[58] = 6'h2b;
        mem[59] = 6'h1f;
        mem[60] = 6'h39;
        mem[61] = 6'h20;
        mem[62] = 6'h17;
        mem[63] = 6'h1c;
    end
endmodule

module odo_sbox_small25(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h00;
        mem[1] = 6'h38;
        mem[2] = 6'h0d;
        mem[3] = 6'h07;
        mem[4] = 6'h0e;
        mem[5] = 6'h2b;
        mem[6] = 6'h33;
        mem[7] = 6'h15;
        mem[8] = 6'h04;
        mem[9] = 6'h2c;
        mem[10] = 6'h13;
        mem[11] = 6'h2d;
        mem[12] = 6'h3e;
        mem[13] = 6'h36;
        mem[14] = 6'h31;
        mem[15] = 6'h05;
        mem[16] = 6'h16;
        mem[17] = 6'h37;
        mem[18] = 6'h1a;
        mem[19] = 6'h25;
        mem[20] = 6'h1d;
        mem[21] = 6'h23;
        mem[22] = 6'h08;
        mem[23] = 6'h3a;
        mem[24] = 6'h0a;
        mem[25] = 6'h35;
        mem[26] = 6'h2e;
        mem[27] = 6'h1c;
        mem[28] = 6'h29;
        mem[29] = 6'h17;
        mem[30] = 6'h26;
        mem[31] = 6'h1b;
        mem[32] = 6'h03;
        mem[33] = 6'h10;
        mem[34] = 6'h1e;
        mem[35] = 6'h2a;
        mem[36] = 6'h14;
        mem[37] = 6'h21;
        mem[38] = 6'h2f;
        mem[39] = 6'h01;
        mem[40] = 6'h30;
        mem[41] = 6'h3b;
        mem[42] = 6'h24;
        mem[43] = 6'h18;
        mem[44] = 6'h0f;
        mem[45] = 6'h3f;
        mem[46] = 6'h27;
        mem[47] = 6'h06;
        mem[48] = 6'h11;
        mem[49] = 6'h09;
        mem[50] = 6'h0c;
        mem[51] = 6'h34;
        mem[52] = 6'h20;
        mem[53] = 6'h12;
        mem[54] = 6'h0b;
        mem[55] = 6'h1f;
        mem[56] = 6'h3d;
        mem[57] = 6'h22;
        mem[58] = 6'h3c;
        mem[59] = 6'h28;
        mem[60] = 6'h39;
        mem[61] = 6'h02;
        mem[62] = 6'h32;
        mem[63] = 6'h19;
    end
endmodule

module odo_sbox_small26(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h34;
        mem[1] = 6'h2f;
        mem[2] = 6'h0d;
        mem[3] = 6'h1d;
        mem[4] = 6'h13;
        mem[5] = 6'h37;
        mem[6] = 6'h2c;
        mem[7] = 6'h1b;
        mem[8] = 6'h0e;
        mem[9] = 6'h03;
        mem[10] = 6'h15;
        mem[11] = 6'h29;
        mem[12] = 6'h35;
        mem[13] = 6'h24;
        mem[14] = 6'h3f;
        mem[15] = 6'h1c;
        mem[16] = 6'h2a;
        mem[17] = 6'h25;
        mem[18] = 6'h1e;
        mem[19] = 6'h01;
        mem[20] = 6'h26;
        mem[21] = 6'h2d;
        mem[22] = 6'h27;
        mem[23] = 6'h0f;
        mem[24] = 6'h3b;
        mem[25] = 6'h2e;
        mem[26] = 6'h28;
        mem[27] = 6'h16;
        mem[28] = 6'h1f;
        mem[29] = 6'h1a;
        mem[30] = 6'h05;
        mem[31] = 6'h12;
        mem[32] = 6'h11;
        mem[33] = 6'h23;
        mem[34] = 6'h20;
        mem[35] = 6'h09;
        mem[36] = 6'h06;
        mem[37] = 6'h0b;
        mem[38] = 6'h18;
        mem[39] = 6'h30;
        mem[40] = 6'h0c;
        mem[41] = 6'h08;
        mem[42] = 6'h32;
        mem[43] = 6'h0a;
        mem[44] = 6'h36;
        mem[45] = 6'h21;
        mem[46] = 6'h00;
        mem[47] = 6'h14;
        mem[48] = 6'h38;
        mem[49] = 6'h31;
        mem[50] = 6'h10;
        mem[51] = 6'h3e;
        mem[52] = 6'h33;
        mem[53] = 6'h19;
        mem[54] = 6'h3d;
        mem[55] = 6'h17;
        mem[56] = 6'h3a;
        mem[57] = 6'h02;
        mem[58] = 6'h07;
        mem[59] = 6'h2b;
        mem[60] = 6'h39;
        mem[61] = 6'h3c;
        mem[62] = 6'h22;
        mem[63] = 6'h04;
    end
endmodule

module odo_sbox_small27(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0b;
        mem[1] = 6'h11;
        mem[2] = 6'h26;
        mem[3] = 6'h25;
        mem[4] = 6'h1e;
        mem[5] = 6'h14;
        mem[6] = 6'h35;
        mem[7] = 6'h32;
        mem[8] = 6'h29;
        mem[9] = 6'h33;
        mem[10] = 6'h3c;
        mem[11] = 6'h0e;
        mem[12] = 6'h24;
        mem[13] = 6'h05;
        mem[14] = 6'h06;
        mem[15] = 6'h39;
        mem[16] = 6'h21;
        mem[17] = 6'h31;
        mem[18] = 6'h2a;
        mem[19] = 6'h1c;
        mem[20] = 6'h3e;
        mem[21] = 6'h2f;
        mem[22] = 6'h36;
        mem[23] = 6'h27;
        mem[24] = 6'h34;
        mem[25] = 6'h1b;
        mem[26] = 6'h0c;
        mem[27] = 6'h04;
        mem[28] = 6'h0f;
        mem[29] = 6'h02;
        mem[30] = 6'h2b;
        mem[31] = 6'h3f;
        mem[32] = 6'h38;
        mem[33] = 6'h30;
        mem[34] = 6'h2d;
        mem[35] = 6'h18;
        mem[36] = 6'h3d;
        mem[37] = 6'h3b;
        mem[38] = 6'h1f;
        mem[39] = 6'h3a;
        mem[40] = 6'h17;
        mem[41] = 6'h10;
        mem[42] = 6'h08;
        mem[43] = 6'h20;
        mem[44] = 6'h09;
        mem[45] = 6'h1a;
        mem[46] = 6'h28;
        mem[47] = 6'h2e;
        mem[48] = 6'h37;
        mem[49] = 6'h00;
        mem[50] = 6'h0d;
        mem[51] = 6'h15;
        mem[52] = 6'h2c;
        mem[53] = 6'h13;
        mem[54] = 6'h01;
        mem[55] = 6'h07;
        mem[56] = 6'h03;
        mem[57] = 6'h16;
        mem[58] = 6'h22;
        mem[59] = 6'h0a;
        mem[60] = 6'h23;
        mem[61] = 6'h19;
        mem[62] = 6'h1d;
        mem[63] = 6'h12;
    end
endmodule

module odo_sbox_small28(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h29;
        mem[1] = 6'h18;
        mem[2] = 6'h17;
        mem[3] = 6'h0c;
        mem[4] = 6'h39;
        mem[5] = 6'h04;
        mem[6] = 6'h0a;
        mem[7] = 6'h25;
        mem[8] = 6'h0e;
        mem[9] = 6'h01;
        mem[10] = 6'h31;
        mem[11] = 6'h1d;
        mem[12] = 6'h22;
        mem[13] = 6'h3c;
        mem[14] = 6'h10;
        mem[15] = 6'h3e;
        mem[16] = 6'h3b;
        mem[17] = 6'h1a;
        mem[18] = 6'h08;
        mem[19] = 6'h37;
        mem[20] = 6'h1e;
        mem[21] = 6'h2e;
        mem[22] = 6'h34;
        mem[23] = 6'h20;
        mem[24] = 6'h2f;
        mem[25] = 6'h32;
        mem[26] = 6'h1f;
        mem[27] = 6'h11;
        mem[28] = 6'h15;
        mem[29] = 6'h35;
        mem[30] = 6'h06;
        mem[31] = 6'h07;
        mem[32] = 6'h2a;
        mem[33] = 6'h02;
        mem[34] = 6'h14;
        mem[35] = 6'h16;
        mem[36] = 6'h00;
        mem[37] = 6'h3d;
        mem[38] = 6'h23;
        mem[39] = 6'h27;
        mem[40] = 6'h0b;
        mem[41] = 6'h28;
        mem[42] = 6'h3a;
        mem[43] = 6'h2c;
        mem[44] = 6'h13;
        mem[45] = 6'h1c;
        mem[46] = 6'h3f;
        mem[47] = 6'h12;
        mem[48] = 6'h03;
        mem[49] = 6'h2d;
        mem[50] = 6'h26;
        mem[51] = 6'h19;
        mem[52] = 6'h21;
        mem[53] = 6'h05;
        mem[54] = 6'h2b;
        mem[55] = 6'h36;
        mem[56] = 6'h1b;
        mem[57] = 6'h38;
        mem[58] = 6'h0d;
        mem[59] = 6'h24;
        mem[60] = 6'h30;
        mem[61] = 6'h0f;
        mem[62] = 6'h09;
        mem[63] = 6'h33;
    end
endmodule

module odo_sbox_small29(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h21;
        mem[1] = 6'h00;
        mem[2] = 6'h0e;
        mem[3] = 6'h2d;
        mem[4] = 6'h33;
        mem[5] = 6'h20;
        mem[6] = 6'h25;
        mem[7] = 6'h2c;
        mem[8] = 6'h1e;
        mem[9] = 6'h1c;
        mem[10] = 6'h08;
        mem[11] = 6'h16;
        mem[12] = 6'h0b;
        mem[13] = 6'h3f;
        mem[14] = 6'h34;
        mem[15] = 6'h35;
        mem[16] = 6'h1f;
        mem[17] = 6'h24;
        mem[18] = 6'h32;
        mem[19] = 6'h2e;
        mem[20] = 6'h19;
        mem[21] = 6'h14;
        mem[22] = 6'h0f;
        mem[23] = 6'h06;
        mem[24] = 6'h2f;
        mem[25] = 6'h39;
        mem[26] = 6'h38;
        mem[27] = 6'h37;
        mem[28] = 6'h0c;
        mem[29] = 6'h13;
        mem[30] = 6'h0a;
        mem[31] = 6'h03;
        mem[32] = 6'h01;
        mem[33] = 6'h02;
        mem[34] = 6'h31;
        mem[35] = 6'h27;
        mem[36] = 6'h23;
        mem[37] = 6'h1b;
        mem[38] = 6'h11;
        mem[39] = 6'h0d;
        mem[40] = 6'h3a;
        mem[41] = 6'h05;
        mem[42] = 6'h15;
        mem[43] = 6'h36;
        mem[44] = 6'h17;
        mem[45] = 6'h10;
        mem[46] = 6'h07;
        mem[47] = 6'h26;
        mem[48] = 6'h3c;
        mem[49] = 6'h09;
        mem[50] = 6'h04;
        mem[51] = 6'h29;
        mem[52] = 6'h1d;
        mem[53] = 6'h12;
        mem[54] = 6'h1a;
        mem[55] = 6'h2b;
        mem[56] = 6'h3b;
        mem[57] = 6'h3d;
        mem[58] = 6'h30;
        mem[59] = 6'h22;
        mem[60] = 6'h2a;
        mem[61] = 6'h18;
        mem[62] = 6'h3e;
        mem[63] = 6'h28;
    end
endmodule

module odo_sbox_small30(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1f;
        mem[1] = 6'h1b;
        mem[2] = 6'h01;
        mem[3] = 6'h11;
        mem[4] = 6'h1a;
        mem[5] = 6'h19;
        mem[6] = 6'h31;
        mem[7] = 6'h07;
        mem[8] = 6'h09;
        mem[9] = 6'h0b;
        mem[10] = 6'h17;
        mem[11] = 6'h08;
        mem[12] = 6'h30;
        mem[13] = 6'h13;
        mem[14] = 6'h3d;
        mem[15] = 6'h2f;
        mem[16] = 6'h1e;
        mem[17] = 6'h04;
        mem[18] = 6'h25;
        mem[19] = 6'h2b;
        mem[20] = 6'h10;
        mem[21] = 6'h12;
        mem[22] = 6'h0d;
        mem[23] = 6'h35;
        mem[24] = 6'h3e;
        mem[25] = 6'h0f;
        mem[26] = 6'h22;
        mem[27] = 6'h05;
        mem[28] = 6'h3f;
        mem[29] = 6'h2a;
        mem[30] = 6'h0c;
        mem[31] = 6'h20;
        mem[32] = 6'h23;
        mem[33] = 6'h32;
        mem[34] = 6'h06;
        mem[35] = 6'h03;
        mem[36] = 6'h2c;
        mem[37] = 6'h36;
        mem[38] = 6'h14;
        mem[39] = 6'h02;
        mem[40] = 6'h18;
        mem[41] = 6'h29;
        mem[42] = 6'h24;
        mem[43] = 6'h3c;
        mem[44] = 6'h00;
        mem[45] = 6'h21;
        mem[46] = 6'h34;
        mem[47] = 6'h15;
        mem[48] = 6'h0a;
        mem[49] = 6'h0e;
        mem[50] = 6'h28;
        mem[51] = 6'h39;
        mem[52] = 6'h3b;
        mem[53] = 6'h3a;
        mem[54] = 6'h2d;
        mem[55] = 6'h1d;
        mem[56] = 6'h2e;
        mem[57] = 6'h33;
        mem[58] = 6'h26;
        mem[59] = 6'h38;
        mem[60] = 6'h37;
        mem[61] = 6'h1c;
        mem[62] = 6'h27;
        mem[63] = 6'h16;
    end
endmodule

module odo_sbox_small31(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h33;
        mem[1] = 6'h1e;
        mem[2] = 6'h11;
        mem[3] = 6'h3d;
        mem[4] = 6'h02;
        mem[5] = 6'h2c;
        mem[6] = 6'h13;
        mem[7] = 6'h07;
        mem[8] = 6'h38;
        mem[9] = 6'h36;
        mem[10] = 6'h0e;
        mem[11] = 6'h12;
        mem[12] = 6'h35;
        mem[13] = 6'h0c;
        mem[14] = 6'h37;
        mem[15] = 6'h31;
        mem[16] = 6'h08;
        mem[17] = 6'h16;
        mem[18] = 6'h05;
        mem[19] = 6'h3a;
        mem[20] = 6'h0f;
        mem[21] = 6'h1f;
        mem[22] = 6'h3f;
        mem[23] = 6'h04;
        mem[24] = 6'h29;
        mem[25] = 6'h15;
        mem[26] = 6'h34;
        mem[27] = 6'h0a;
        mem[28] = 6'h19;
        mem[29] = 6'h2b;
        mem[30] = 6'h32;
        mem[31] = 6'h00;
        mem[32] = 6'h3b;
        mem[33] = 6'h21;
        mem[34] = 6'h2a;
        mem[35] = 6'h0b;
        mem[36] = 6'h20;
        mem[37] = 6'h24;
        mem[38] = 6'h17;
        mem[39] = 6'h09;
        mem[40] = 6'h39;
        mem[41] = 6'h14;
        mem[42] = 6'h27;
        mem[43] = 6'h06;
        mem[44] = 6'h3e;
        mem[45] = 6'h18;
        mem[46] = 6'h0d;
        mem[47] = 6'h23;
        mem[48] = 6'h22;
        mem[49] = 6'h01;
        mem[50] = 6'h1a;
        mem[51] = 6'h1b;
        mem[52] = 6'h3c;
        mem[53] = 6'h26;
        mem[54] = 6'h10;
        mem[55] = 6'h2e;
        mem[56] = 6'h1c;
        mem[57] = 6'h30;
        mem[58] = 6'h2d;
        mem[59] = 6'h25;
        mem[60] = 6'h03;
        mem[61] = 6'h28;
        mem[62] = 6'h2f;
        mem[63] = 6'h1d;
    end
endmodule

module odo_sbox_small32(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h13;
        mem[1] = 6'h18;
        mem[2] = 6'h37;
        mem[3] = 6'h1f;
        mem[4] = 6'h10;
        mem[5] = 6'h02;
        mem[6] = 6'h07;
        mem[7] = 6'h28;
        mem[8] = 6'h21;
        mem[9] = 6'h16;
        mem[10] = 6'h34;
        mem[11] = 6'h0b;
        mem[12] = 6'h2c;
        mem[13] = 6'h0d;
        mem[14] = 6'h17;
        mem[15] = 6'h0f;
        mem[16] = 6'h11;
        mem[17] = 6'h25;
        mem[18] = 6'h15;
        mem[19] = 6'h1e;
        mem[20] = 6'h3c;
        mem[21] = 6'h2e;
        mem[22] = 6'h35;
        mem[23] = 6'h29;
        mem[24] = 6'h05;
        mem[25] = 6'h0e;
        mem[26] = 6'h06;
        mem[27] = 6'h1a;
        mem[28] = 6'h1c;
        mem[29] = 6'h3f;
        mem[30] = 6'h03;
        mem[31] = 6'h31;
        mem[32] = 6'h0a;
        mem[33] = 6'h27;
        mem[34] = 6'h36;
        mem[35] = 6'h26;
        mem[36] = 6'h39;
        mem[37] = 6'h19;
        mem[38] = 6'h24;
        mem[39] = 6'h00;
        mem[40] = 6'h2d;
        mem[41] = 6'h3a;
        mem[42] = 6'h2f;
        mem[43] = 6'h08;
        mem[44] = 6'h33;
        mem[45] = 6'h3e;
        mem[46] = 6'h2a;
        mem[47] = 6'h1b;
        mem[48] = 6'h30;
        mem[49] = 6'h32;
        mem[50] = 6'h12;
        mem[51] = 6'h14;
        mem[52] = 6'h22;
        mem[53] = 6'h1d;
        mem[54] = 6'h09;
        mem[55] = 6'h0c;
        mem[56] = 6'h01;
        mem[57] = 6'h23;
        mem[58] = 6'h3b;
        mem[59] = 6'h38;
        mem[60] = 6'h20;
        mem[61] = 6'h2b;
        mem[62] = 6'h04;
        mem[63] = 6'h3d;
    end
endmodule

module odo_sbox_small33(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h31;
        mem[1] = 6'h1b;
        mem[2] = 6'h24;
        mem[3] = 6'h11;
        mem[4] = 6'h10;
        mem[5] = 6'h3a;
        mem[6] = 6'h26;
        mem[7] = 6'h1a;
        mem[8] = 6'h1e;
        mem[9] = 6'h1d;
        mem[10] = 6'h22;
        mem[11] = 6'h17;
        mem[12] = 6'h0c;
        mem[13] = 6'h19;
        mem[14] = 6'h16;
        mem[15] = 6'h3c;
        mem[16] = 6'h0f;
        mem[17] = 6'h35;
        mem[18] = 6'h12;
        mem[19] = 6'h30;
        mem[20] = 6'h39;
        mem[21] = 6'h2e;
        mem[22] = 6'h27;
        mem[23] = 6'h28;
        mem[24] = 6'h08;
        mem[25] = 6'h0e;
        mem[26] = 6'h21;
        mem[27] = 6'h2a;
        mem[28] = 6'h2d;
        mem[29] = 6'h23;
        mem[30] = 6'h3e;
        mem[31] = 6'h07;
        mem[32] = 6'h25;
        mem[33] = 6'h13;
        mem[34] = 6'h36;
        mem[35] = 6'h0a;
        mem[36] = 6'h3d;
        mem[37] = 6'h15;
        mem[38] = 6'h0d;
        mem[39] = 6'h14;
        mem[40] = 6'h34;
        mem[41] = 6'h09;
        mem[42] = 6'h2b;
        mem[43] = 6'h3b;
        mem[44] = 6'h1f;
        mem[45] = 6'h03;
        mem[46] = 6'h2c;
        mem[47] = 6'h05;
        mem[48] = 6'h01;
        mem[49] = 6'h29;
        mem[50] = 6'h02;
        mem[51] = 6'h2f;
        mem[52] = 6'h37;
        mem[53] = 6'h18;
        mem[54] = 6'h00;
        mem[55] = 6'h38;
        mem[56] = 6'h04;
        mem[57] = 6'h20;
        mem[58] = 6'h3f;
        mem[59] = 6'h06;
        mem[60] = 6'h33;
        mem[61] = 6'h1c;
        mem[62] = 6'h0b;
        mem[63] = 6'h32;
    end
endmodule

module odo_sbox_small34(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h39;
        mem[1] = 6'h23;
        mem[2] = 6'h1e;
        mem[3] = 6'h13;
        mem[4] = 6'h2d;
        mem[5] = 6'h10;
        mem[6] = 6'h26;
        mem[7] = 6'h07;
        mem[8] = 6'h3c;
        mem[9] = 6'h0e;
        mem[10] = 6'h1c;
        mem[11] = 6'h17;
        mem[12] = 6'h2c;
        mem[13] = 6'h30;
        mem[14] = 6'h04;
        mem[15] = 6'h11;
        mem[16] = 6'h37;
        mem[17] = 6'h0a;
        mem[18] = 6'h2a;
        mem[19] = 6'h1f;
        mem[20] = 6'h0b;
        mem[21] = 6'h21;
        mem[22] = 6'h0f;
        mem[23] = 6'h3a;
        mem[24] = 6'h0d;
        mem[25] = 6'h32;
        mem[26] = 6'h0c;
        mem[27] = 6'h34;
        mem[28] = 6'h25;
        mem[29] = 6'h09;
        mem[30] = 6'h3b;
        mem[31] = 6'h24;
        mem[32] = 6'h31;
        mem[33] = 6'h35;
        mem[34] = 6'h00;
        mem[35] = 6'h3e;
        mem[36] = 6'h1d;
        mem[37] = 6'h1a;
        mem[38] = 6'h03;
        mem[39] = 6'h08;
        mem[40] = 6'h27;
        mem[41] = 6'h2e;
        mem[42] = 6'h02;
        mem[43] = 6'h3d;
        mem[44] = 6'h38;
        mem[45] = 6'h01;
        mem[46] = 6'h18;
        mem[47] = 6'h3f;
        mem[48] = 6'h1b;
        mem[49] = 6'h36;
        mem[50] = 6'h29;
        mem[51] = 6'h06;
        mem[52] = 6'h19;
        mem[53] = 6'h12;
        mem[54] = 6'h22;
        mem[55] = 6'h2f;
        mem[56] = 6'h15;
        mem[57] = 6'h20;
        mem[58] = 6'h2b;
        mem[59] = 6'h33;
        mem[60] = 6'h05;
        mem[61] = 6'h28;
        mem[62] = 6'h14;
        mem[63] = 6'h16;
    end
endmodule

module odo_sbox_small35(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0d;
        mem[1] = 6'h08;
        mem[2] = 6'h2b;
        mem[3] = 6'h1a;
        mem[4] = 6'h2f;
        mem[5] = 6'h32;
        mem[6] = 6'h39;
        mem[7] = 6'h1c;
        mem[8] = 6'h03;
        mem[9] = 6'h13;
        mem[10] = 6'h00;
        mem[11] = 6'h1f;
        mem[12] = 6'h3b;
        mem[13] = 6'h31;
        mem[14] = 6'h01;
        mem[15] = 6'h22;
        mem[16] = 6'h09;
        mem[17] = 6'h06;
        mem[18] = 6'h34;
        mem[19] = 6'h19;
        mem[20] = 6'h16;
        mem[21] = 6'h3f;
        mem[22] = 6'h27;
        mem[23] = 6'h14;
        mem[24] = 6'h3d;
        mem[25] = 6'h35;
        mem[26] = 6'h38;
        mem[27] = 6'h3a;
        mem[28] = 6'h18;
        mem[29] = 6'h24;
        mem[30] = 6'h25;
        mem[31] = 6'h2c;
        mem[32] = 6'h2d;
        mem[33] = 6'h0e;
        mem[34] = 6'h3e;
        mem[35] = 6'h0f;
        mem[36] = 6'h0c;
        mem[37] = 6'h28;
        mem[38] = 6'h0b;
        mem[39] = 6'h30;
        mem[40] = 6'h29;
        mem[41] = 6'h2a;
        mem[42] = 6'h10;
        mem[43] = 6'h1b;
        mem[44] = 6'h36;
        mem[45] = 6'h11;
        mem[46] = 6'h04;
        mem[47] = 6'h15;
        mem[48] = 6'h21;
        mem[49] = 6'h02;
        mem[50] = 6'h07;
        mem[51] = 6'h37;
        mem[52] = 6'h23;
        mem[53] = 6'h33;
        mem[54] = 6'h0a;
        mem[55] = 6'h2e;
        mem[56] = 6'h05;
        mem[57] = 6'h20;
        mem[58] = 6'h1d;
        mem[59] = 6'h26;
        mem[60] = 6'h17;
        mem[61] = 6'h3c;
        mem[62] = 6'h12;
        mem[63] = 6'h1e;
    end
endmodule

module odo_sbox_small36(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h22;
        mem[1] = 6'h2c;
        mem[2] = 6'h1e;
        mem[3] = 6'h0c;
        mem[4] = 6'h29;
        mem[5] = 6'h28;
        mem[6] = 6'h18;
        mem[7] = 6'h11;
        mem[8] = 6'h03;
        mem[9] = 6'h1b;
        mem[10] = 6'h13;
        mem[11] = 6'h0f;
        mem[12] = 6'h2e;
        mem[13] = 6'h2f;
        mem[14] = 6'h2a;
        mem[15] = 6'h12;
        mem[16] = 6'h20;
        mem[17] = 6'h23;
        mem[18] = 6'h38;
        mem[19] = 6'h26;
        mem[20] = 6'h3c;
        mem[21] = 6'h04;
        mem[22] = 6'h33;
        mem[23] = 6'h35;
        mem[24] = 6'h0a;
        mem[25] = 6'h3b;
        mem[26] = 6'h05;
        mem[27] = 6'h21;
        mem[28] = 6'h3d;
        mem[29] = 6'h1f;
        mem[30] = 6'h00;
        mem[31] = 6'h2b;
        mem[32] = 6'h0d;
        mem[33] = 6'h16;
        mem[34] = 6'h1d;
        mem[35] = 6'h0b;
        mem[36] = 6'h32;
        mem[37] = 6'h30;
        mem[38] = 6'h17;
        mem[39] = 6'h08;
        mem[40] = 6'h3e;
        mem[41] = 6'h39;
        mem[42] = 6'h07;
        mem[43] = 6'h31;
        mem[44] = 6'h1a;
        mem[45] = 6'h25;
        mem[46] = 6'h1c;
        mem[47] = 6'h15;
        mem[48] = 6'h02;
        mem[49] = 6'h24;
        mem[50] = 6'h01;
        mem[51] = 6'h10;
        mem[52] = 6'h2d;
        mem[53] = 6'h06;
        mem[54] = 6'h27;
        mem[55] = 6'h09;
        mem[56] = 6'h34;
        mem[57] = 6'h36;
        mem[58] = 6'h14;
        mem[59] = 6'h19;
        mem[60] = 6'h3f;
        mem[61] = 6'h3a;
        mem[62] = 6'h0e;
        mem[63] = 6'h37;
    end
endmodule

module odo_sbox_small37(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h17;
        mem[1] = 6'h10;
        mem[2] = 6'h2b;
        mem[3] = 6'h12;
        mem[4] = 6'h3e;
        mem[5] = 6'h02;
        mem[6] = 6'h33;
        mem[7] = 6'h3c;
        mem[8] = 6'h13;
        mem[9] = 6'h06;
        mem[10] = 6'h31;
        mem[11] = 6'h2c;
        mem[12] = 6'h3f;
        mem[13] = 6'h09;
        mem[14] = 6'h34;
        mem[15] = 6'h01;
        mem[16] = 6'h05;
        mem[17] = 6'h0e;
        mem[18] = 6'h1b;
        mem[19] = 6'h1f;
        mem[20] = 6'h26;
        mem[21] = 6'h30;
        mem[22] = 6'h36;
        mem[23] = 6'h00;
        mem[24] = 6'h11;
        mem[25] = 6'h3b;
        mem[26] = 6'h38;
        mem[27] = 6'h07;
        mem[28] = 6'h18;
        mem[29] = 6'h0b;
        mem[30] = 6'h3d;
        mem[31] = 6'h1a;
        mem[32] = 6'h08;
        mem[33] = 6'h03;
        mem[34] = 6'h39;
        mem[35] = 6'h2e;
        mem[36] = 6'h1e;
        mem[37] = 6'h21;
        mem[38] = 6'h22;
        mem[39] = 6'h19;
        mem[40] = 6'h32;
        mem[41] = 6'h2f;
        mem[42] = 6'h2d;
        mem[43] = 6'h0a;
        mem[44] = 6'h16;
        mem[45] = 6'h15;
        mem[46] = 6'h28;
        mem[47] = 6'h0f;
        mem[48] = 6'h1d;
        mem[49] = 6'h37;
        mem[50] = 6'h29;
        mem[51] = 6'h23;
        mem[52] = 6'h2a;
        mem[53] = 6'h1c;
        mem[54] = 6'h0c;
        mem[55] = 6'h14;
        mem[56] = 6'h27;
        mem[57] = 6'h25;
        mem[58] = 6'h04;
        mem[59] = 6'h20;
        mem[60] = 6'h0d;
        mem[61] = 6'h35;
        mem[62] = 6'h24;
        mem[63] = 6'h3a;
    end
endmodule

module odo_sbox_small38(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h14;
        mem[1] = 6'h09;
        mem[2] = 6'h37;
        mem[3] = 6'h1c;
        mem[4] = 6'h15;
        mem[5] = 6'h03;
        mem[6] = 6'h12;
        mem[7] = 6'h35;
        mem[8] = 6'h2e;
        mem[9] = 6'h18;
        mem[10] = 6'h30;
        mem[11] = 6'h1e;
        mem[12] = 6'h3f;
        mem[13] = 6'h00;
        mem[14] = 6'h3c;
        mem[15] = 6'h23;
        mem[16] = 6'h31;
        mem[17] = 6'h1f;
        mem[18] = 6'h06;
        mem[19] = 6'h08;
        mem[20] = 6'h16;
        mem[21] = 6'h27;
        mem[22] = 6'h36;
        mem[23] = 6'h19;
        mem[24] = 6'h25;
        mem[25] = 6'h2b;
        mem[26] = 6'h02;
        mem[27] = 6'h10;
        mem[28] = 6'h22;
        mem[29] = 6'h2a;
        mem[30] = 6'h39;
        mem[31] = 6'h0c;
        mem[32] = 6'h05;
        mem[33] = 6'h1d;
        mem[34] = 6'h38;
        mem[35] = 6'h17;
        mem[36] = 6'h33;
        mem[37] = 6'h0b;
        mem[38] = 6'h1a;
        mem[39] = 6'h29;
        mem[40] = 6'h3b;
        mem[41] = 6'h07;
        mem[42] = 6'h20;
        mem[43] = 6'h2f;
        mem[44] = 6'h21;
        mem[45] = 6'h28;
        mem[46] = 6'h32;
        mem[47] = 6'h26;
        mem[48] = 6'h0e;
        mem[49] = 6'h3a;
        mem[50] = 6'h13;
        mem[51] = 6'h2c;
        mem[52] = 6'h01;
        mem[53] = 6'h04;
        mem[54] = 6'h1b;
        mem[55] = 6'h34;
        mem[56] = 6'h11;
        mem[57] = 6'h3e;
        mem[58] = 6'h24;
        mem[59] = 6'h0f;
        mem[60] = 6'h3d;
        mem[61] = 6'h2d;
        mem[62] = 6'h0d;
        mem[63] = 6'h0a;
    end
endmodule

module odo_sbox_small39(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h26;
        mem[1] = 6'h3d;
        mem[2] = 6'h1e;
        mem[3] = 6'h3c;
        mem[4] = 6'h12;
        mem[5] = 6'h2a;
        mem[6] = 6'h33;
        mem[7] = 6'h0a;
        mem[8] = 6'h25;
        mem[9] = 6'h2d;
        mem[10] = 6'h14;
        mem[11] = 6'h20;
        mem[12] = 6'h24;
        mem[13] = 6'h2b;
        mem[14] = 6'h0d;
        mem[15] = 6'h27;
        mem[16] = 6'h06;
        mem[17] = 6'h23;
        mem[18] = 6'h29;
        mem[19] = 6'h09;
        mem[20] = 6'h31;
        mem[21] = 6'h36;
        mem[22] = 6'h22;
        mem[23] = 6'h17;
        mem[24] = 6'h30;
        mem[25] = 6'h2f;
        mem[26] = 6'h1d;
        mem[27] = 6'h08;
        mem[28] = 6'h05;
        mem[29] = 6'h32;
        mem[30] = 6'h0c;
        mem[31] = 6'h11;
        mem[32] = 6'h2c;
        mem[33] = 6'h1c;
        mem[34] = 6'h34;
        mem[35] = 6'h02;
        mem[36] = 6'h0f;
        mem[37] = 6'h18;
        mem[38] = 6'h2e;
        mem[39] = 6'h1f;
        mem[40] = 6'h38;
        mem[41] = 6'h04;
        mem[42] = 6'h35;
        mem[43] = 6'h15;
        mem[44] = 6'h3f;
        mem[45] = 6'h0b;
        mem[46] = 6'h3a;
        mem[47] = 6'h28;
        mem[48] = 6'h07;
        mem[49] = 6'h13;
        mem[50] = 6'h00;
        mem[51] = 6'h3b;
        mem[52] = 6'h39;
        mem[53] = 6'h37;
        mem[54] = 6'h03;
        mem[55] = 6'h19;
        mem[56] = 6'h3e;
        mem[57] = 6'h10;
        mem[58] = 6'h1b;
        mem[59] = 6'h16;
        mem[60] = 6'h01;
        mem[61] = 6'h21;
        mem[62] = 6'h1a;
        mem[63] = 6'h0e;
    end
endmodule

module odo_sbox_large0(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h174;
        mem[1] = 10'h089;
        mem[2] = 10'h108;
        mem[3] = 10'h3a0;
        mem[4] = 10'h1c7;
        mem[5] = 10'h0f3;
        mem[6] = 10'h3a7;
        mem[7] = 10'h05a;
        mem[8] = 10'h181;
        mem[9] = 10'h3b3;
        mem[10] = 10'h0ee;
        mem[11] = 10'h3f0;
        mem[12] = 10'h299;
        mem[13] = 10'h1a9;
        mem[14] = 10'h0f7;
        mem[15] = 10'h378;
        mem[16] = 10'h0f8;
        mem[17] = 10'h0a9;
        mem[18] = 10'h3c7;
        mem[19] = 10'h3f9;
        mem[20] = 10'h385;
        mem[21] = 10'h118;
        mem[22] = 10'h1dc;
        mem[23] = 10'h333;
        mem[24] = 10'h32f;
        mem[25] = 10'h04c;
        mem[26] = 10'h3eb;
        mem[27] = 10'h1b4;
        mem[28] = 10'h1ff;
        mem[29] = 10'h38b;
        mem[30] = 10'h3de;
        mem[31] = 10'h3b2;
        mem[32] = 10'h1f1;
        mem[33] = 10'h0d6;
        mem[34] = 10'h001;
        mem[35] = 10'h2bd;
        mem[36] = 10'h353;
        mem[37] = 10'h067;
        mem[38] = 10'h31f;
        mem[39] = 10'h3a5;
        mem[40] = 10'h2ae;
        mem[41] = 10'h0a7;
        mem[42] = 10'h222;
        mem[43] = 10'h101;
        mem[44] = 10'h317;
        mem[45] = 10'h1c6;
        mem[46] = 10'h37c;
        mem[47] = 10'h2f0;
        mem[48] = 10'h26f;
        mem[49] = 10'h30b;
        mem[50] = 10'h207;
        mem[51] = 10'h08b;
        mem[52] = 10'h21f;
        mem[53] = 10'h17b;
        mem[54] = 10'h0cc;
        mem[55] = 10'h136;
        mem[56] = 10'h096;
        mem[57] = 10'h3ea;
        mem[58] = 10'h0b0;
        mem[59] = 10'h052;
        mem[60] = 10'h03d;
        mem[61] = 10'h2ce;
        mem[62] = 10'h252;
        mem[63] = 10'h07c;
        mem[64] = 10'h1c0;
        mem[65] = 10'h006;
        mem[66] = 10'h19a;
        mem[67] = 10'h33f;
        mem[68] = 10'h0c0;
        mem[69] = 10'h1b3;
        mem[70] = 10'h1d4;
        mem[71] = 10'h0e6;
        mem[72] = 10'h0c8;
        mem[73] = 10'h20a;
        mem[74] = 10'h30f;
        mem[75] = 10'h2e2;
        mem[76] = 10'h397;
        mem[77] = 10'h0d7;
        mem[78] = 10'h1c3;
        mem[79] = 10'h330;
        mem[80] = 10'h3fb;
        mem[81] = 10'h226;
        mem[82] = 10'h2dc;
        mem[83] = 10'h3b1;
        mem[84] = 10'h0c7;
        mem[85] = 10'h3e1;
        mem[86] = 10'h1f3;
        mem[87] = 10'h0fa;
        mem[88] = 10'h2e1;
        mem[89] = 10'h0d5;
        mem[90] = 10'h0a5;
        mem[91] = 10'h371;
        mem[92] = 10'h112;
        mem[93] = 10'h39b;
        mem[94] = 10'h34e;
        mem[95] = 10'h0fd;
        mem[96] = 10'h3ee;
        mem[97] = 10'h042;
        mem[98] = 10'h216;
        mem[99] = 10'h314;
        mem[100] = 10'h139;
        mem[101] = 10'h2d9;
        mem[102] = 10'h018;
        mem[103] = 10'h06c;
        mem[104] = 10'h0c4;
        mem[105] = 10'h0e4;
        mem[106] = 10'h37f;
        mem[107] = 10'h2c8;
        mem[108] = 10'h1cf;
        mem[109] = 10'h3fe;
        mem[110] = 10'h1b5;
        mem[111] = 10'h256;
        mem[112] = 10'h1ca;
        mem[113] = 10'h1dd;
        mem[114] = 10'h0d3;
        mem[115] = 10'h223;
        mem[116] = 10'h260;
        mem[117] = 10'h295;
        mem[118] = 10'h3b0;
        mem[119] = 10'h110;
        mem[120] = 10'h12c;
        mem[121] = 10'h28b;
        mem[122] = 10'h0fb;
        mem[123] = 10'h0ea;
        mem[124] = 10'h220;
        mem[125] = 10'h2c6;
        mem[126] = 10'h3f4;
        mem[127] = 10'h19f;
        mem[128] = 10'h01f;
        mem[129] = 10'h19c;
        mem[130] = 10'h1d2;
        mem[131] = 10'h153;
        mem[132] = 10'h233;
        mem[133] = 10'h1e3;
        mem[134] = 10'h094;
        mem[135] = 10'h24b;
        mem[136] = 10'h321;
        mem[137] = 10'h2b0;
        mem[138] = 10'h305;
        mem[139] = 10'h08a;
        mem[140] = 10'h0cd;
        mem[141] = 10'h2e6;
        mem[142] = 10'h0f0;
        mem[143] = 10'h2fe;
        mem[144] = 10'h1fb;
        mem[145] = 10'h13f;
        mem[146] = 10'h3ca;
        mem[147] = 10'h278;
        mem[148] = 10'h360;
        mem[149] = 10'h248;
        mem[150] = 10'h064;
        mem[151] = 10'h0fe;
        mem[152] = 10'h1c9;
        mem[153] = 10'h092;
        mem[154] = 10'h365;
        mem[155] = 10'h1d1;
        mem[156] = 10'h24e;
        mem[157] = 10'h085;
        mem[158] = 10'h28f;
        mem[159] = 10'h1a8;
        mem[160] = 10'h281;
        mem[161] = 10'h356;
        mem[162] = 10'h057;
        mem[163] = 10'h3ba;
        mem[164] = 10'h106;
        mem[165] = 10'h218;
        mem[166] = 10'h17f;
        mem[167] = 10'h2d6;
        mem[168] = 10'h104;
        mem[169] = 10'h351;
        mem[170] = 10'h190;
        mem[171] = 10'h1f0;
        mem[172] = 10'h189;
        mem[173] = 10'h120;
        mem[174] = 10'h099;
        mem[175] = 10'h1a6;
        mem[176] = 10'h277;
        mem[177] = 10'h3ed;
        mem[178] = 10'h045;
        mem[179] = 10'h3e4;
        mem[180] = 10'h39c;
        mem[181] = 10'h38d;
        mem[182] = 10'h33e;
        mem[183] = 10'h023;
        mem[184] = 10'h06f;
        mem[185] = 10'h1df;
        mem[186] = 10'h381;
        mem[187] = 10'h1a3;
        mem[188] = 10'h255;
        mem[189] = 10'h0f2;
        mem[190] = 10'h3d9;
        mem[191] = 10'h362;
        mem[192] = 10'h3d1;
        mem[193] = 10'h066;
        mem[194] = 10'h11c;
        mem[195] = 10'h322;
        mem[196] = 10'h2d4;
        mem[197] = 10'h152;
        mem[198] = 10'h114;
        mem[199] = 10'h199;
        mem[200] = 10'h291;
        mem[201] = 10'h228;
        mem[202] = 10'h34f;
        mem[203] = 10'h399;
        mem[204] = 10'h1a5;
        mem[205] = 10'h079;
        mem[206] = 10'h249;
        mem[207] = 10'h0d2;
        mem[208] = 10'h168;
        mem[209] = 10'h2cd;
        mem[210] = 10'h0e3;
        mem[211] = 10'h225;
        mem[212] = 10'h1db;
        mem[213] = 10'h03b;
        mem[214] = 10'h350;
        mem[215] = 10'h18c;
        mem[216] = 10'h14c;
        mem[217] = 10'h27b;
        mem[218] = 10'h032;
        mem[219] = 10'h01d;
        mem[220] = 10'h352;
        mem[221] = 10'h2c9;
        mem[222] = 10'h185;
        mem[223] = 10'h2e3;
        mem[224] = 10'h021;
        mem[225] = 10'h2ba;
        mem[226] = 10'h176;
        mem[227] = 10'h020;
        mem[228] = 10'h320;
        mem[229] = 10'h19b;
        mem[230] = 10'h326;
        mem[231] = 10'h076;
        mem[232] = 10'h323;
        mem[233] = 10'h221;
        mem[234] = 10'h366;
        mem[235] = 10'h3d5;
        mem[236] = 10'h2a1;
        mem[237] = 10'h25c;
        mem[238] = 10'h00c;
        mem[239] = 10'h15f;
        mem[240] = 10'h270;
        mem[241] = 10'h227;
        mem[242] = 10'h2ab;
        mem[243] = 10'h003;
        mem[244] = 10'h375;
        mem[245] = 10'h318;
        mem[246] = 10'h05c;
        mem[247] = 10'h0bf;
        mem[248] = 10'h16e;
        mem[249] = 10'h2da;
        mem[250] = 10'h15a;
        mem[251] = 10'h17c;
        mem[252] = 10'h387;
        mem[253] = 10'h103;
        mem[254] = 10'h049;
        mem[255] = 10'h29e;
        mem[256] = 10'h05e;
        mem[257] = 10'h027;
        mem[258] = 10'h135;
        mem[259] = 10'h04f;
        mem[260] = 10'h11f;
        mem[261] = 10'h20f;
        mem[262] = 10'h034;
        mem[263] = 10'h395;
        mem[264] = 10'h148;
        mem[265] = 10'h20d;
        mem[266] = 10'h008;
        mem[267] = 10'h23b;
        mem[268] = 10'h2e9;
        mem[269] = 10'h327;
        mem[270] = 10'h048;
        mem[271] = 10'h1ee;
        mem[272] = 10'h18b;
        mem[273] = 10'h398;
        mem[274] = 10'h07d;
        mem[275] = 10'h3ac;
        mem[276] = 10'h259;
        mem[277] = 10'h2be;
        mem[278] = 10'h025;
        mem[279] = 10'h00e;
        mem[280] = 10'h02d;
        mem[281] = 10'h1c8;
        mem[282] = 10'h175;
        mem[283] = 10'h211;
        mem[284] = 10'h364;
        mem[285] = 10'h344;
        mem[286] = 10'h06e;
        mem[287] = 10'h328;
        mem[288] = 10'h0af;
        mem[289] = 10'h24d;
        mem[290] = 10'h1fe;
        mem[291] = 10'h1b6;
        mem[292] = 10'h3ef;
        mem[293] = 10'h28e;
        mem[294] = 10'h2f2;
        mem[295] = 10'h23e;
        mem[296] = 10'h232;
        mem[297] = 10'h0f4;
        mem[298] = 10'h290;
        mem[299] = 10'h279;
        mem[300] = 10'h1d3;
        mem[301] = 10'h15c;
        mem[302] = 10'h131;
        mem[303] = 10'h1ef;
        mem[304] = 10'h037;
        mem[305] = 10'h16b;
        mem[306] = 10'h3a2;
        mem[307] = 10'h3a8;
        mem[308] = 10'h15e;
        mem[309] = 10'h21e;
        mem[310] = 10'h3ff;
        mem[311] = 10'h186;
        mem[312] = 10'h38c;
        mem[313] = 10'h149;
        mem[314] = 10'h3ce;
        mem[315] = 10'h22c;
        mem[316] = 10'h2c0;
        mem[317] = 10'h14e;
        mem[318] = 10'h164;
        mem[319] = 10'h235;
        mem[320] = 10'h111;
        mem[321] = 10'h3a4;
        mem[322] = 10'h029;
        mem[323] = 10'h293;
        mem[324] = 10'h17d;
        mem[325] = 10'h31e;
        mem[326] = 10'h22b;
        mem[327] = 10'h03e;
        mem[328] = 10'h1cc;
        mem[329] = 10'h010;
        mem[330] = 10'h004;
        mem[331] = 10'h0b2;
        mem[332] = 10'h3c6;
        mem[333] = 10'h179;
        mem[334] = 10'h1e2;
        mem[335] = 10'h083;
        mem[336] = 10'h10a;
        mem[337] = 10'h144;
        mem[338] = 10'h240;
        mem[339] = 10'h288;
        mem[340] = 10'h055;
        mem[341] = 10'h0d1;
        mem[342] = 10'h147;
        mem[343] = 10'h126;
        mem[344] = 10'h1af;
        mem[345] = 10'h391;
        mem[346] = 10'h347;
        mem[347] = 10'h1f9;
        mem[348] = 10'h1c2;
        mem[349] = 10'h3d4;
        mem[350] = 10'h08e;
        mem[351] = 10'h196;
        mem[352] = 10'h332;
        mem[353] = 10'h25e;
        mem[354] = 10'h3c1;
        mem[355] = 10'h35f;
        mem[356] = 10'h158;
        mem[357] = 10'h0ad;
        mem[358] = 10'h0db;
        mem[359] = 10'h0a0;
        mem[360] = 10'h033;
        mem[361] = 10'h204;
        mem[362] = 10'h05b;
        mem[363] = 10'h07b;
        mem[364] = 10'h23d;
        mem[365] = 10'h1a0;
        mem[366] = 10'h22f;
        mem[367] = 10'h34b;
        mem[368] = 10'h1cd;
        mem[369] = 10'h2a7;
        mem[370] = 10'h33b;
        mem[371] = 10'h271;
        mem[372] = 10'h246;
        mem[373] = 10'h11e;
        mem[374] = 10'h3c0;
        mem[375] = 10'h081;
        mem[376] = 10'h234;
        mem[377] = 10'h2b8;
        mem[378] = 10'h369;
        mem[379] = 10'h251;
        mem[380] = 10'h146;
        mem[381] = 10'h262;
        mem[382] = 10'h302;
        mem[383] = 10'h348;
        mem[384] = 10'h2cf;
        mem[385] = 10'h261;
        mem[386] = 10'h123;
        mem[387] = 10'h3cc;
        mem[388] = 10'h1cb;
        mem[389] = 10'h12f;
        mem[390] = 10'h29b;
        mem[391] = 10'h1e9;
        mem[392] = 10'h264;
        mem[393] = 10'h016;
        mem[394] = 10'h0ca;
        mem[395] = 10'h2a3;
        mem[396] = 10'h1ba;
        mem[397] = 10'h05f;
        mem[398] = 10'h041;
        mem[399] = 10'h184;
        mem[400] = 10'h343;
        mem[401] = 10'h14b;
        mem[402] = 10'h340;
        mem[403] = 10'h337;
        mem[404] = 10'h0b3;
        mem[405] = 10'h265;
        mem[406] = 10'h2b6;
        mem[407] = 10'h368;
        mem[408] = 10'h0ba;
        mem[409] = 10'h0e7;
        mem[410] = 10'h070;
        mem[411] = 10'h253;
        mem[412] = 10'h028;
        mem[413] = 10'h3c3;
        mem[414] = 10'h39f;
        mem[415] = 10'h0ed;
        mem[416] = 10'h090;
        mem[417] = 10'h1a1;
        mem[418] = 10'h27e;
        mem[419] = 10'h31d;
        mem[420] = 10'h0bc;
        mem[421] = 10'h200;
        mem[422] = 10'h354;
        mem[423] = 10'h1b0;
        mem[424] = 10'h019;
        mem[425] = 10'h237;
        mem[426] = 10'h2b7;
        mem[427] = 10'h053;
        mem[428] = 10'h134;
        mem[429] = 10'h289;
        mem[430] = 10'h38e;
        mem[431] = 10'h014;
        mem[432] = 10'h21c;
        mem[433] = 10'h062;
        mem[434] = 10'h312;
        mem[435] = 10'h3ae;
        mem[436] = 10'h1ab;
        mem[437] = 10'h115;
        mem[438] = 10'h043;
        mem[439] = 10'h121;
        mem[440] = 10'h0e0;
        mem[441] = 10'h0ce;
        mem[442] = 10'h017;
        mem[443] = 10'h3e2;
        mem[444] = 10'h238;
        mem[445] = 10'h357;
        mem[446] = 10'h14f;
        mem[447] = 10'h1f6;
        mem[448] = 10'h250;
        mem[449] = 10'h074;
        mem[450] = 10'h0c6;
        mem[451] = 10'h180;
        mem[452] = 10'h379;
        mem[453] = 10'h0cf;
        mem[454] = 10'h26d;
        mem[455] = 10'h2a4;
        mem[456] = 10'h283;
        mem[457] = 10'h159;
        mem[458] = 10'h269;
        mem[459] = 10'h0d0;
        mem[460] = 10'h268;
        mem[461] = 10'h36e;
        mem[462] = 10'h2eb;
        mem[463] = 10'h3bb;
        mem[464] = 10'h39e;
        mem[465] = 10'h3da;
        mem[466] = 10'h031;
        mem[467] = 10'h1da;
        mem[468] = 10'h298;
        mem[469] = 10'h2e5;
        mem[470] = 10'h33d;
        mem[471] = 10'h372;
        mem[472] = 10'h292;
        mem[473] = 10'h063;
        mem[474] = 10'h2b9;
        mem[475] = 10'h358;
        mem[476] = 10'h0df;
        mem[477] = 10'h0fc;
        mem[478] = 10'h35b;
        mem[479] = 10'h32a;
        mem[480] = 10'h214;
        mem[481] = 10'h2d8;
        mem[482] = 10'h308;
        mem[483] = 10'h0c1;
        mem[484] = 10'h306;
        mem[485] = 10'h191;
        mem[486] = 10'h307;
        mem[487] = 10'h3d6;
        mem[488] = 10'h217;
        mem[489] = 10'h17a;
        mem[490] = 10'h3e6;
        mem[491] = 10'h282;
        mem[492] = 10'h3d8;
        mem[493] = 10'h338;
        mem[494] = 10'h0b8;
        mem[495] = 10'h1bf;
        mem[496] = 10'h3f8;
        mem[497] = 10'h009;
        mem[498] = 10'h37d;
        mem[499] = 10'h384;
        mem[500] = 10'h087;
        mem[501] = 10'h0a1;
        mem[502] = 10'h3e8;
        mem[503] = 10'h241;
        mem[504] = 10'h022;
        mem[505] = 10'h3cb;
        mem[506] = 10'h1fa;
        mem[507] = 10'h16d;
        mem[508] = 10'h39d;
        mem[509] = 10'h08f;
        mem[510] = 10'h16c;
        mem[511] = 10'h155;
        mem[512] = 10'h061;
        mem[513] = 10'h22a;
        mem[514] = 10'h3f2;
        mem[515] = 10'h0f9;
        mem[516] = 10'h396;
        mem[517] = 10'h005;
        mem[518] = 10'h3db;
        mem[519] = 10'h236;
        mem[520] = 10'h2ad;
        mem[521] = 10'h361;
        mem[522] = 10'h2a5;
        mem[523] = 10'h1fc;
        mem[524] = 10'h2d5;
        mem[525] = 10'h00f;
        mem[526] = 10'h07f;
        mem[527] = 10'h35d;
        mem[528] = 10'h2ef;
        mem[529] = 10'h09a;
        mem[530] = 10'h209;
        mem[531] = 10'h142;
        mem[532] = 10'h0b4;
        mem[533] = 10'h1d9;
        mem[534] = 10'h26b;
        mem[535] = 10'h138;
        mem[536] = 10'h331;
        mem[537] = 10'h20c;
        mem[538] = 10'h160;
        mem[539] = 10'h27c;
        mem[540] = 10'h2aa;
        mem[541] = 10'h208;
        mem[542] = 10'h18a;
        mem[543] = 10'h09b;
        mem[544] = 10'h21a;
        mem[545] = 10'h00b;
        mem[546] = 10'h097;
        mem[547] = 10'h34a;
        mem[548] = 10'h32b;
        mem[549] = 10'h000;
        mem[550] = 10'h301;
        mem[551] = 10'h215;
        mem[552] = 10'h377;
        mem[553] = 10'h13d;
        mem[554] = 10'h1bc;
        mem[555] = 10'h01e;
        mem[556] = 10'h355;
        mem[557] = 10'h172;
        mem[558] = 10'h346;
        mem[559] = 10'h1c5;
        mem[560] = 10'h3f3;
        mem[561] = 10'h19d;
        mem[562] = 10'h3fd;
        mem[563] = 10'h3e0;
        mem[564] = 10'h1de;
        mem[565] = 10'h1f4;
        mem[566] = 10'h3ec;
        mem[567] = 10'h0c5;
        mem[568] = 10'h3d0;
        mem[569] = 10'h22d;
        mem[570] = 10'h165;
        mem[571] = 10'h2d1;
        mem[572] = 10'h2f5;
        mem[573] = 10'h1d6;
        mem[574] = 10'h18d;
        mem[575] = 10'h170;
        mem[576] = 10'h210;
        mem[577] = 10'h2bb;
        mem[578] = 10'h2f1;
        mem[579] = 10'h177;
        mem[580] = 10'h2b4;
        mem[581] = 10'h263;
        mem[582] = 10'h124;
        mem[583] = 10'h00d;
        mem[584] = 10'h31b;
        mem[585] = 10'h2c4;
        mem[586] = 10'h266;
        mem[587] = 10'h125;
        mem[588] = 10'h2df;
        mem[589] = 10'h339;
        mem[590] = 10'h082;
        mem[591] = 10'h002;
        mem[592] = 10'h25d;
        mem[593] = 10'h276;
        mem[594] = 10'h224;
        mem[595] = 10'h0b6;
        mem[596] = 10'h015;
        mem[597] = 10'h151;
        mem[598] = 10'h056;
        mem[599] = 10'h192;
        mem[600] = 10'h047;
        mem[601] = 10'h3b4;
        mem[602] = 10'h068;
        mem[603] = 10'h0e5;
        mem[604] = 10'h0e8;
        mem[605] = 10'h194;
        mem[606] = 10'h335;
        mem[607] = 10'h3cd;
        mem[608] = 10'h3f5;
        mem[609] = 10'h13a;
        mem[610] = 10'h3f1;
        mem[611] = 10'h21b;
        mem[612] = 10'h09f;
        mem[613] = 10'h030;
        mem[614] = 10'h14a;
        mem[615] = 10'h28a;
        mem[616] = 10'h119;
        mem[617] = 10'h2a2;
        mem[618] = 10'h35a;
        mem[619] = 10'h05d;
        mem[620] = 10'h3af;
        mem[621] = 10'h128;
        mem[622] = 10'h03f;
        mem[623] = 10'h376;
        mem[624] = 10'h3a9;
        mem[625] = 10'h1bd;
        mem[626] = 10'h20b;
        mem[627] = 10'h245;
        mem[628] = 10'h035;
        mem[629] = 10'h0a2;
        mem[630] = 10'h109;
        mem[631] = 10'h26e;
        mem[632] = 10'h23f;
        mem[633] = 10'h1ce;
        mem[634] = 10'h161;
        mem[635] = 10'h2dd;
        mem[636] = 10'h2ec;
        mem[637] = 10'h2a9;
        mem[638] = 10'h37e;
        mem[639] = 10'h230;
        mem[640] = 10'h01c;
        mem[641] = 10'h145;
        mem[642] = 10'h374;
        mem[643] = 10'h0ab;
        mem[644] = 10'h23a;
        mem[645] = 10'h03c;
        mem[646] = 10'h0dc;
        mem[647] = 10'h206;
        mem[648] = 10'h31c;
        mem[649] = 10'h2cb;
        mem[650] = 10'h26a;
        mem[651] = 10'h162;
        mem[652] = 10'h013;
        mem[653] = 10'h349;
        mem[654] = 10'h3dc;
        mem[655] = 10'h050;
        mem[656] = 10'h0da;
        mem[657] = 10'h257;
        mem[658] = 10'h1d8;
        mem[659] = 10'h32c;
        mem[660] = 10'h2b3;
        mem[661] = 10'h18e;
        mem[662] = 10'h3ad;
        mem[663] = 10'h1f2;
        mem[664] = 10'h1c4;
        mem[665] = 10'h1eb;
        mem[666] = 10'h0ef;
        mem[667] = 10'h0be;
        mem[668] = 10'h3cf;
        mem[669] = 10'h0f5;
        mem[670] = 10'h0f1;
        mem[671] = 10'h1e4;
        mem[672] = 10'h20e;
        mem[673] = 10'h065;
        mem[674] = 10'h09c;
        mem[675] = 10'h116;
        mem[676] = 10'h071;
        mem[677] = 10'h3c2;
        mem[678] = 10'h202;
        mem[679] = 10'h198;
        mem[680] = 10'h28c;
        mem[681] = 10'h163;
        mem[682] = 10'h3df;
        mem[683] = 10'h3fc;
        mem[684] = 10'h02c;
        mem[685] = 10'h19e;
        mem[686] = 10'h2bf;
        mem[687] = 10'h1be;
        mem[688] = 10'h29c;
        mem[689] = 10'h2b5;
        mem[690] = 10'h213;
        mem[691] = 10'h102;
        mem[692] = 10'h32e;
        mem[693] = 10'h09d;
        mem[694] = 10'h2e4;
        mem[695] = 10'h12a;
        mem[696] = 10'h388;
        mem[697] = 10'h0f6;
        mem[698] = 10'h1ed;
        mem[699] = 10'h02b;
        mem[700] = 10'h33a;
        mem[701] = 10'h122;
        mem[702] = 10'h2a8;
        mem[703] = 10'h2d3;
        mem[704] = 10'h1e8;
        mem[705] = 10'h2b2;
        mem[706] = 10'h2db;
        mem[707] = 10'h0aa;
        mem[708] = 10'h093;
        mem[709] = 10'h060;
        mem[710] = 10'h1b2;
        mem[711] = 10'h11d;
        mem[712] = 10'h267;
        mem[713] = 10'h304;
        mem[714] = 10'h34d;
        mem[715] = 10'h036;
        mem[716] = 10'h300;
        mem[717] = 10'h12b;
        mem[718] = 10'h25b;
        mem[719] = 10'h0d9;
        mem[720] = 10'h130;
        mem[721] = 10'h113;
        mem[722] = 10'h150;
        mem[723] = 10'h3e9;
        mem[724] = 10'h100;
        mem[725] = 10'h383;
        mem[726] = 10'h244;
        mem[727] = 10'h078;
        mem[728] = 10'h239;
        mem[729] = 10'h35e;
        mem[730] = 10'h393;
        mem[731] = 10'h1a7;
        mem[732] = 10'h2ee;
        mem[733] = 10'h183;
        mem[734] = 10'h2e8;
        mem[735] = 10'h10c;
        mem[736] = 10'h32d;
        mem[737] = 10'h3a3;
        mem[738] = 10'h2f3;
        mem[739] = 10'h098;
        mem[740] = 10'h0ff;
        mem[741] = 10'h36f;
        mem[742] = 10'h247;
        mem[743] = 10'h2c7;
        mem[744] = 10'h2f7;
        mem[745] = 10'h0b5;
        mem[746] = 10'h3c4;
        mem[747] = 10'h0b1;
        mem[748] = 10'h0a6;
        mem[749] = 10'h02f;
        mem[750] = 10'h143;
        mem[751] = 10'h011;
        mem[752] = 10'h2d7;
        mem[753] = 10'h2c2;
        mem[754] = 10'h0e1;
        mem[755] = 10'h2fd;
        mem[756] = 10'h342;
        mem[757] = 10'h044;
        mem[758] = 10'h205;
        mem[759] = 10'h1a2;
        mem[760] = 10'h334;
        mem[761] = 10'h3d2;
        mem[762] = 10'h095;
        mem[763] = 10'h127;
        mem[764] = 10'h27f;
        mem[765] = 10'h3dd;
        mem[766] = 10'h2e0;
        mem[767] = 10'h367;
        mem[768] = 10'h0cb;
        mem[769] = 10'h3e5;
        mem[770] = 10'h197;
        mem[771] = 10'h12e;
        mem[772] = 10'h1b8;
        mem[773] = 10'h0c2;
        mem[774] = 10'h00a;
        mem[775] = 10'h26c;
        mem[776] = 10'h3d3;
        mem[777] = 10'h07e;
        mem[778] = 10'h0c9;
        mem[779] = 10'h1b7;
        mem[780] = 10'h10b;
        mem[781] = 10'h37b;
        mem[782] = 10'h154;
        mem[783] = 10'h3bf;
        mem[784] = 10'h12d;
        mem[785] = 10'h02a;
        mem[786] = 10'h13b;
        mem[787] = 10'h316;
        mem[788] = 10'h024;
        mem[789] = 10'h3e3;
        mem[790] = 10'h2f6;
        mem[791] = 10'h077;
        mem[792] = 10'h258;
        mem[793] = 10'h394;
        mem[794] = 10'h0ec;
        mem[795] = 10'h3bd;
        mem[796] = 10'h11a;
        mem[797] = 10'h072;
        mem[798] = 10'h1a4;
        mem[799] = 10'h242;
        mem[800] = 10'h1fd;
        mem[801] = 10'h1ae;
        mem[802] = 10'h3c5;
        mem[803] = 10'h30a;
        mem[804] = 10'h311;
        mem[805] = 10'h380;
        mem[806] = 10'h2ea;
        mem[807] = 10'h363;
        mem[808] = 10'h3fa;
        mem[809] = 10'h09e;
        mem[810] = 10'h178;
        mem[811] = 10'h0d8;
        mem[812] = 10'h34c;
        mem[813] = 10'h193;
        mem[814] = 10'h3d7;
        mem[815] = 10'h02e;
        mem[816] = 10'h15b;
        mem[817] = 10'h06b;
        mem[818] = 10'h182;
        mem[819] = 10'h16a;
        mem[820] = 10'h392;
        mem[821] = 10'h166;
        mem[822] = 10'h30e;
        mem[823] = 10'h01b;
        mem[824] = 10'h2c3;
        mem[825] = 10'h046;
        mem[826] = 10'h026;
        mem[827] = 10'h3ab;
        mem[828] = 10'h10f;
        mem[829] = 10'h2cc;
        mem[830] = 10'h286;
        mem[831] = 10'h31a;
        mem[832] = 10'h3b9;
        mem[833] = 10'h1e7;
        mem[834] = 10'h382;
        mem[835] = 10'h294;
        mem[836] = 10'h187;
        mem[837] = 10'h229;
        mem[838] = 10'h36d;
        mem[839] = 10'h07a;
        mem[840] = 10'h132;
        mem[841] = 10'h105;
        mem[842] = 10'h06d;
        mem[843] = 10'h2d0;
        mem[844] = 10'h0bd;
        mem[845] = 10'h080;
        mem[846] = 10'h2a0;
        mem[847] = 10'h273;
        mem[848] = 10'h073;
        mem[849] = 10'h373;
        mem[850] = 10'h390;
        mem[851] = 10'h280;
        mem[852] = 10'h0ae;
        mem[853] = 10'h140;
        mem[854] = 10'h3f7;
        mem[855] = 10'h0de;
        mem[856] = 10'h3a6;
        mem[857] = 10'h133;
        mem[858] = 10'h0a4;
        mem[859] = 10'h2de;
        mem[860] = 10'h171;
        mem[861] = 10'h18f;
        mem[862] = 10'h274;
        mem[863] = 10'h13c;
        mem[864] = 10'h296;
        mem[865] = 10'h2bc;
        mem[866] = 10'h2c1;
        mem[867] = 10'h0d4;
        mem[868] = 10'h059;
        mem[869] = 10'h173;
        mem[870] = 10'h359;
        mem[871] = 10'h039;
        mem[872] = 10'h3be;
        mem[873] = 10'h1b9;
        mem[874] = 10'h086;
        mem[875] = 10'h169;
        mem[876] = 10'h272;
        mem[877] = 10'h06a;
        mem[878] = 10'h051;
        mem[879] = 10'h0e9;
        mem[880] = 10'h22e;
        mem[881] = 10'h007;
        mem[882] = 10'h38f;
        mem[883] = 10'h2ff;
        mem[884] = 10'h08d;
        mem[885] = 10'h17e;
        mem[886] = 10'h29a;
        mem[887] = 10'h284;
        mem[888] = 10'h36b;
        mem[889] = 10'h04a;
        mem[890] = 10'h329;
        mem[891] = 10'h1f5;
        mem[892] = 10'h23c;
        mem[893] = 10'h1e0;
        mem[894] = 10'h1ec;
        mem[895] = 10'h219;
        mem[896] = 10'h370;
        mem[897] = 10'h1d0;
        mem[898] = 10'h29d;
        mem[899] = 10'h325;
        mem[900] = 10'h3c9;
        mem[901] = 10'h0a8;
        mem[902] = 10'h3aa;
        mem[903] = 10'h0bb;
        mem[904] = 10'h341;
        mem[905] = 10'h0a3;
        mem[906] = 10'h012;
        mem[907] = 10'h231;
        mem[908] = 10'h2f8;
        mem[909] = 10'h04d;
        mem[910] = 10'h1c1;
        mem[911] = 10'h054;
        mem[912] = 10'h1d5;
        mem[913] = 10'h15d;
        mem[914] = 10'h2f4;
        mem[915] = 10'h275;
        mem[916] = 10'h3e7;
        mem[917] = 10'h27d;
        mem[918] = 10'h1e6;
        mem[919] = 10'h091;
        mem[920] = 10'h37a;
        mem[921] = 10'h3c8;
        mem[922] = 10'h3a1;
        mem[923] = 10'h157;
        mem[924] = 10'h10d;
        mem[925] = 10'h167;
        mem[926] = 10'h107;
        mem[927] = 10'h2fb;
        mem[928] = 10'h2e7;
        mem[929] = 10'h075;
        mem[930] = 10'h25a;
        mem[931] = 10'h309;
        mem[932] = 10'h2d2;
        mem[933] = 10'h0e2;
        mem[934] = 10'h0ac;
        mem[935] = 10'h0c3;
        mem[936] = 10'h1ad;
        mem[937] = 10'h2fa;
        mem[938] = 10'h03a;
        mem[939] = 10'h01a;
        mem[940] = 10'h2c5;
        mem[941] = 10'h1b1;
        mem[942] = 10'h2ed;
        mem[943] = 10'h310;
        mem[944] = 10'h3b6;
        mem[945] = 10'h1e5;
        mem[946] = 10'h3f6;
        mem[947] = 10'h0b9;
        mem[948] = 10'h3b7;
        mem[949] = 10'h203;
        mem[950] = 10'h285;
        mem[951] = 10'h13e;
        mem[952] = 10'h39a;
        mem[953] = 10'h36a;
        mem[954] = 10'h129;
        mem[955] = 10'h315;
        mem[956] = 10'h3bc;
        mem[957] = 10'h038;
        mem[958] = 10'h30c;
        mem[959] = 10'h24c;
        mem[960] = 10'h38a;
        mem[961] = 10'h29f;
        mem[962] = 10'h2f9;
        mem[963] = 10'h35c;
        mem[964] = 10'h137;
        mem[965] = 10'h04e;
        mem[966] = 10'h088;
        mem[967] = 10'h3b5;
        mem[968] = 10'h2ac;
        mem[969] = 10'h389;
        mem[970] = 10'h30d;
        mem[971] = 10'h2fc;
        mem[972] = 10'h2b1;
        mem[973] = 10'h16f;
        mem[974] = 10'h2ca;
        mem[975] = 10'h141;
        mem[976] = 10'h0eb;
        mem[977] = 10'h28d;
        mem[978] = 10'h1d7;
        mem[979] = 10'h336;
        mem[980] = 10'h254;
        mem[981] = 10'h21d;
        mem[982] = 10'h04b;
        mem[983] = 10'h084;
        mem[984] = 10'h386;
        mem[985] = 10'h2a6;
        mem[986] = 10'h117;
        mem[987] = 10'h24a;
        mem[988] = 10'h319;
        mem[989] = 10'h2af;
        mem[990] = 10'h1bb;
        mem[991] = 10'h297;
        mem[992] = 10'h36c;
        mem[993] = 10'h212;
        mem[994] = 10'h14d;
        mem[995] = 10'h201;
        mem[996] = 10'h345;
        mem[997] = 10'h0dd;
        mem[998] = 10'h10e;
        mem[999] = 10'h313;
        mem[1000] = 10'h1e1;
        mem[1001] = 10'h1f7;
        mem[1002] = 10'h1ac;
        mem[1003] = 10'h156;
        mem[1004] = 10'h1ea;
        mem[1005] = 10'h08c;
        mem[1006] = 10'h069;
        mem[1007] = 10'h24f;
        mem[1008] = 10'h324;
        mem[1009] = 10'h33c;
        mem[1010] = 10'h303;
        mem[1011] = 10'h1aa;
        mem[1012] = 10'h195;
        mem[1013] = 10'h243;
        mem[1014] = 10'h058;
        mem[1015] = 10'h040;
        mem[1016] = 10'h0b7;
        mem[1017] = 10'h11b;
        mem[1018] = 10'h287;
        mem[1019] = 10'h27a;
        mem[1020] = 10'h188;
        mem[1021] = 10'h1f8;
        mem[1022] = 10'h3b8;
        mem[1023] = 10'h25f;
    end
endmodule

module odo_sbox_large1(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h0c3;
        mem[1] = 10'h18b;
        mem[2] = 10'h1e4;
        mem[3] = 10'h081;
        mem[4] = 10'h123;
        mem[5] = 10'h095;
        mem[6] = 10'h107;
        mem[7] = 10'h229;
        mem[8] = 10'h3fc;
        mem[9] = 10'h225;
        mem[10] = 10'h125;
        mem[11] = 10'h388;
        mem[12] = 10'h266;
        mem[13] = 10'h291;
        mem[14] = 10'h1df;
        mem[15] = 10'h0cd;
        mem[16] = 10'h31a;
        mem[17] = 10'h0dd;
        mem[18] = 10'h167;
        mem[19] = 10'h284;
        mem[20] = 10'h27c;
        mem[21] = 10'h271;
        mem[22] = 10'h041;
        mem[23] = 10'h398;
        mem[24] = 10'h36a;
        mem[25] = 10'h0c4;
        mem[26] = 10'h108;
        mem[27] = 10'h272;
        mem[28] = 10'h042;
        mem[29] = 10'h3b8;
        mem[30] = 10'h08b;
        mem[31] = 10'h317;
        mem[32] = 10'h013;
        mem[33] = 10'h1b8;
        mem[34] = 10'h0fb;
        mem[35] = 10'h03e;
        mem[36] = 10'h176;
        mem[37] = 10'h2e2;
        mem[38] = 10'h1cd;
        mem[39] = 10'h394;
        mem[40] = 10'h0f6;
        mem[41] = 10'h39b;
        mem[42] = 10'h0c6;
        mem[43] = 10'h06f;
        mem[44] = 10'h3a6;
        mem[45] = 10'h1b7;
        mem[46] = 10'h189;
        mem[47] = 10'h355;
        mem[48] = 10'h14c;
        mem[49] = 10'h0d4;
        mem[50] = 10'h024;
        mem[51] = 10'h21c;
        mem[52] = 10'h0a9;
        mem[53] = 10'h227;
        mem[54] = 10'h142;
        mem[55] = 10'h019;
        mem[56] = 10'h2b3;
        mem[57] = 10'h0e9;
        mem[58] = 10'h3f4;
        mem[59] = 10'h1e3;
        mem[60] = 10'h1f1;
        mem[61] = 10'h11b;
        mem[62] = 10'h2ab;
        mem[63] = 10'h34e;
        mem[64] = 10'h2a8;
        mem[65] = 10'h0b0;
        mem[66] = 10'h131;
        mem[67] = 10'h078;
        mem[68] = 10'h2fe;
        mem[69] = 10'h0e4;
        mem[70] = 10'h001;
        mem[71] = 10'h2fd;
        mem[72] = 10'h141;
        mem[73] = 10'h3de;
        mem[74] = 10'h1c1;
        mem[75] = 10'h19f;
        mem[76] = 10'h285;
        mem[77] = 10'h187;
        mem[78] = 10'h279;
        mem[79] = 10'h1b6;
        mem[80] = 10'h339;
        mem[81] = 10'h15e;
        mem[82] = 10'h055;
        mem[83] = 10'h08f;
        mem[84] = 10'h37d;
        mem[85] = 10'h114;
        mem[86] = 10'h216;
        mem[87] = 10'h1cf;
        mem[88] = 10'h36c;
        mem[89] = 10'h02e;
        mem[90] = 10'h274;
        mem[91] = 10'h19e;
        mem[92] = 10'h0b6;
        mem[93] = 10'h133;
        mem[94] = 10'h07a;
        mem[95] = 10'h166;
        mem[96] = 10'h038;
        mem[97] = 10'h3c5;
        mem[98] = 10'h3b0;
        mem[99] = 10'h180;
        mem[100] = 10'h14b;
        mem[101] = 10'h061;
        mem[102] = 10'h380;
        mem[103] = 10'h09a;
        mem[104] = 10'h3bb;
        mem[105] = 10'h391;
        mem[106] = 10'h080;
        mem[107] = 10'h260;
        mem[108] = 10'h3df;
        mem[109] = 10'h3e5;
        mem[110] = 10'h359;
        mem[111] = 10'h0f7;
        mem[112] = 10'h2f5;
        mem[113] = 10'h2c7;
        mem[114] = 10'h16c;
        mem[115] = 10'h002;
        mem[116] = 10'h022;
        mem[117] = 10'h3fb;
        mem[118] = 10'h35b;
        mem[119] = 10'h2b8;
        mem[120] = 10'h105;
        mem[121] = 10'h033;
        mem[122] = 10'h0c2;
        mem[123] = 10'h22f;
        mem[124] = 10'h164;
        mem[125] = 10'h3fe;
        mem[126] = 10'h344;
        mem[127] = 10'h1da;
        mem[128] = 10'h008;
        mem[129] = 10'h157;
        mem[130] = 10'h3d0;
        mem[131] = 10'h3a7;
        mem[132] = 10'h1c0;
        mem[133] = 10'h28c;
        mem[134] = 10'h162;
        mem[135] = 10'h09c;
        mem[136] = 10'h38f;
        mem[137] = 10'h3e8;
        mem[138] = 10'h1ef;
        mem[139] = 10'h25b;
        mem[140] = 10'h32e;
        mem[141] = 10'h202;
        mem[142] = 10'h336;
        mem[143] = 10'h19c;
        mem[144] = 10'h2b4;
        mem[145] = 10'h348;
        mem[146] = 10'h2c1;
        mem[147] = 10'h262;
        mem[148] = 10'h1f3;
        mem[149] = 10'h0d0;
        mem[150] = 10'h2c2;
        mem[151] = 10'h2b1;
        mem[152] = 10'h39e;
        mem[153] = 10'h3b5;
        mem[154] = 10'h315;
        mem[155] = 10'h2fc;
        mem[156] = 10'h383;
        mem[157] = 10'h342;
        mem[158] = 10'h1db;
        mem[159] = 10'h13a;
        mem[160] = 10'h352;
        mem[161] = 10'h1be;
        mem[162] = 10'h1ce;
        mem[163] = 10'h2b9;
        mem[164] = 10'h0ea;
        mem[165] = 10'h2df;
        mem[166] = 10'h045;
        mem[167] = 10'h137;
        mem[168] = 10'h151;
        mem[169] = 10'h34c;
        mem[170] = 10'h3b6;
        mem[171] = 10'h26f;
        mem[172] = 10'h2de;
        mem[173] = 10'h26e;
        mem[174] = 10'h1c8;
        mem[175] = 10'h390;
        mem[176] = 10'h0e6;
        mem[177] = 10'h07c;
        mem[178] = 10'h350;
        mem[179] = 10'h1b2;
        mem[180] = 10'h244;
        mem[181] = 10'h28d;
        mem[182] = 10'h3d5;
        mem[183] = 10'h2f4;
        mem[184] = 10'h124;
        mem[185] = 10'h149;
        mem[186] = 10'h0fd;
        mem[187] = 10'h12d;
        mem[188] = 10'h0f4;
        mem[189] = 10'h27d;
        mem[190] = 10'h33e;
        mem[191] = 10'h31e;
        mem[192] = 10'h302;
        mem[193] = 10'h35c;
        mem[194] = 10'h0ee;
        mem[195] = 10'h313;
        mem[196] = 10'h12c;
        mem[197] = 10'h2db;
        mem[198] = 10'h2f8;
        mem[199] = 10'h08a;
        mem[200] = 10'h2a2;
        mem[201] = 10'h368;
        mem[202] = 10'h395;
        mem[203] = 10'h12b;
        mem[204] = 10'h32f;
        mem[205] = 10'h307;
        mem[206] = 10'h14f;
        mem[207] = 10'h23e;
        mem[208] = 10'h2e1;
        mem[209] = 10'h21a;
        mem[210] = 10'h1fb;
        mem[211] = 10'h258;
        mem[212] = 10'h1b9;
        mem[213] = 10'h0da;
        mem[214] = 10'h33f;
        mem[215] = 10'h268;
        mem[216] = 10'h1fd;
        mem[217] = 10'h059;
        mem[218] = 10'h24a;
        mem[219] = 10'h1ee;
        mem[220] = 10'h292;
        mem[221] = 10'h1f0;
        mem[222] = 10'h1c6;
        mem[223] = 10'h2c8;
        mem[224] = 10'h0a3;
        mem[225] = 10'h161;
        mem[226] = 10'h029;
        mem[227] = 10'h24d;
        mem[228] = 10'h11d;
        mem[229] = 10'h208;
        mem[230] = 10'h2c0;
        mem[231] = 10'h2e3;
        mem[232] = 10'h2d2;
        mem[233] = 10'h06e;
        mem[234] = 10'h090;
        mem[235] = 10'h058;
        mem[236] = 10'h060;
        mem[237] = 10'h231;
        mem[238] = 10'h2b7;
        mem[239] = 10'h1c9;
        mem[240] = 10'h1a8;
        mem[241] = 10'h34f;
        mem[242] = 10'h28f;
        mem[243] = 10'h1b4;
        mem[244] = 10'h26b;
        mem[245] = 10'h386;
        mem[246] = 10'h000;
        mem[247] = 10'h1e8;
        mem[248] = 10'h01d;
        mem[249] = 10'h064;
        mem[250] = 10'h035;
        mem[251] = 10'h286;
        mem[252] = 10'h3cc;
        mem[253] = 10'h147;
        mem[254] = 10'h3ac;
        mem[255] = 10'h102;
        mem[256] = 10'h09b;
        mem[257] = 10'h2af;
        mem[258] = 10'h1d2;
        mem[259] = 10'h299;
        mem[260] = 10'h201;
        mem[261] = 10'h11f;
        mem[262] = 10'h067;
        mem[263] = 10'h053;
        mem[264] = 10'h205;
        mem[265] = 10'h22b;
        mem[266] = 10'h213;
        mem[267] = 10'h121;
        mem[268] = 10'h36e;
        mem[269] = 10'h329;
        mem[270] = 10'h0c9;
        mem[271] = 10'h3d7;
        mem[272] = 10'h016;
        mem[273] = 10'h17f;
        mem[274] = 10'h0a6;
        mem[275] = 10'h1bc;
        mem[276] = 10'h297;
        mem[277] = 10'h35a;
        mem[278] = 10'h10b;
        mem[279] = 10'h3b7;
        mem[280] = 10'h209;
        mem[281] = 10'h075;
        mem[282] = 10'h3ec;
        mem[283] = 10'h2ad;
        mem[284] = 10'h106;
        mem[285] = 10'h24c;
        mem[286] = 10'h1dd;
        mem[287] = 10'h1cc;
        mem[288] = 10'h3c3;
        mem[289] = 10'h0a2;
        mem[290] = 10'h301;
        mem[291] = 10'h369;
        mem[292] = 10'h276;
        mem[293] = 10'h294;
        mem[294] = 10'h2be;
        mem[295] = 10'h1c4;
        mem[296] = 10'h2d1;
        mem[297] = 10'h159;
        mem[298] = 10'h0ff;
        mem[299] = 10'h331;
        mem[300] = 10'h377;
        mem[301] = 10'h278;
        mem[302] = 10'h293;
        mem[303] = 10'h257;
        mem[304] = 10'h3aa;
        mem[305] = 10'h3cb;
        mem[306] = 10'h109;
        mem[307] = 10'h1ad;
        mem[308] = 10'h3b2;
        mem[309] = 10'h117;
        mem[310] = 10'h347;
        mem[311] = 10'h158;
        mem[312] = 10'h2cb;
        mem[313] = 10'h308;
        mem[314] = 10'h044;
        mem[315] = 10'h223;
        mem[316] = 10'h38e;
        mem[317] = 10'h1a1;
        mem[318] = 10'h046;
        mem[319] = 10'h039;
        mem[320] = 10'h1f7;
        mem[321] = 10'h0df;
        mem[322] = 10'h093;
        mem[323] = 10'h20f;
        mem[324] = 10'h06c;
        mem[325] = 10'h305;
        mem[326] = 10'h3c9;
        mem[327] = 10'h30b;
        mem[328] = 10'h22e;
        mem[329] = 10'h13d;
        mem[330] = 10'h296;
        mem[331] = 10'h310;
        mem[332] = 10'h0d7;
        mem[333] = 10'h312;
        mem[334] = 10'h111;
        mem[335] = 10'h140;
        mem[336] = 10'h007;
        mem[337] = 10'h006;
        mem[338] = 10'h13f;
        mem[339] = 10'h0de;
        mem[340] = 10'h207;
        mem[341] = 10'h256;
        mem[342] = 10'h21f;
        mem[343] = 10'h119;
        mem[344] = 10'h0db;
        mem[345] = 10'h0d2;
        mem[346] = 10'h251;
        mem[347] = 10'h054;
        mem[348] = 10'h2f0;
        mem[349] = 10'h2a0;
        mem[350] = 10'h2ee;
        mem[351] = 10'h037;
        mem[352] = 10'h063;
        mem[353] = 10'h0ce;
        mem[354] = 10'h1e6;
        mem[355] = 10'h04a;
        mem[356] = 10'h1c5;
        mem[357] = 10'h2a4;
        mem[358] = 10'h212;
        mem[359] = 10'h238;
        mem[360] = 10'h26a;
        mem[361] = 10'h1ea;
        mem[362] = 10'h387;
        mem[363] = 10'h330;
        mem[364] = 10'h26c;
        mem[365] = 10'h195;
        mem[366] = 10'h1eb;
        mem[367] = 10'h3cd;
        mem[368] = 10'h2e0;
        mem[369] = 10'h3f8;
        mem[370] = 10'h152;
        mem[371] = 10'h017;
        mem[372] = 10'h3d9;
        mem[373] = 10'h2eb;
        mem[374] = 10'h077;
        mem[375] = 10'h37e;
        mem[376] = 10'h03b;
        mem[377] = 10'h1d5;
        mem[378] = 10'h0e8;
        mem[379] = 10'h3d2;
        mem[380] = 10'h071;
        mem[381] = 10'h052;
        mem[382] = 10'h3a9;
        mem[383] = 10'h0c8;
        mem[384] = 10'h25a;
        mem[385] = 10'h217;
        mem[386] = 10'h199;
        mem[387] = 10'h0ac;
        mem[388] = 10'h11c;
        mem[389] = 10'h00b;
        mem[390] = 10'h18c;
        mem[391] = 10'h31f;
        mem[392] = 10'h3b3;
        mem[393] = 10'h19b;
        mem[394] = 10'h0b5;
        mem[395] = 10'h129;
        mem[396] = 10'h1b0;
        mem[397] = 10'h1a5;
        mem[398] = 10'h110;
        mem[399] = 10'h18f;
        mem[400] = 10'h20b;
        mem[401] = 10'h00c;
        mem[402] = 10'h3a4;
        mem[403] = 10'h29b;
        mem[404] = 10'h049;
        mem[405] = 10'h0ca;
        mem[406] = 10'h3e4;
        mem[407] = 10'h3c6;
        mem[408] = 10'h0ae;
        mem[409] = 10'h3e3;
        mem[410] = 10'h0f9;
        mem[411] = 10'h245;
        mem[412] = 10'h0e7;
        mem[413] = 10'h120;
        mem[414] = 10'h05e;
        mem[415] = 10'h24e;
        mem[416] = 10'h204;
        mem[417] = 10'h1ab;
        mem[418] = 10'h335;
        mem[419] = 10'h337;
        mem[420] = 10'h242;
        mem[421] = 10'h1af;
        mem[422] = 10'h0f1;
        mem[423] = 10'h29c;
        mem[424] = 10'h333;
        mem[425] = 10'h15a;
        mem[426] = 10'h39d;
        mem[427] = 10'h236;
        mem[428] = 10'h0ed;
        mem[429] = 10'h08d;
        mem[430] = 10'h115;
        mem[431] = 10'h21e;
        mem[432] = 10'h27f;
        mem[433] = 10'h372;
        mem[434] = 10'h353;
        mem[435] = 10'h02d;
        mem[436] = 10'h215;
        mem[437] = 10'h0c7;
        mem[438] = 10'h364;
        mem[439] = 10'h2b6;
        mem[440] = 10'h0a4;
        mem[441] = 10'h057;
        mem[442] = 10'h22a;
        mem[443] = 10'h254;
        mem[444] = 10'h0a0;
        mem[445] = 10'h1a3;
        mem[446] = 10'h16a;
        mem[447] = 10'h03f;
        mem[448] = 10'h349;
        mem[449] = 10'h338;
        mem[450] = 10'h3fa;
        mem[451] = 10'h39c;
        mem[452] = 10'h3fd;
        mem[453] = 10'h263;
        mem[454] = 10'h28b;
        mem[455] = 10'h0cf;
        mem[456] = 10'h0c5;
        mem[457] = 10'h321;
        mem[458] = 10'h182;
        mem[459] = 10'h3ab;
        mem[460] = 10'h1b1;
        mem[461] = 10'h343;
        mem[462] = 10'h089;
        mem[463] = 10'h2fb;
        mem[464] = 10'h306;
        mem[465] = 10'h1e2;
        mem[466] = 10'h31b;
        mem[467] = 10'h1e0;
        mem[468] = 10'h156;
        mem[469] = 10'h30c;
        mem[470] = 10'h32a;
        mem[471] = 10'h05b;
        mem[472] = 10'h1ac;
        mem[473] = 10'h3e1;
        mem[474] = 10'h17d;
        mem[475] = 10'h2a9;
        mem[476] = 10'h32d;
        mem[477] = 10'h134;
        mem[478] = 10'h2cf;
        mem[479] = 10'h2e8;
        mem[480] = 10'h088;
        mem[481] = 10'h191;
        mem[482] = 10'h1a2;
        mem[483] = 10'h094;
        mem[484] = 10'h08c;
        mem[485] = 10'h051;
        mem[486] = 10'h309;
        mem[487] = 10'h3f0;
        mem[488] = 10'h0b1;
        mem[489] = 10'h0ab;
        mem[490] = 10'h3c7;
        mem[491] = 10'h37c;
        mem[492] = 10'h085;
        mem[493] = 10'h10c;
        mem[494] = 10'h340;
        mem[495] = 10'h050;
        mem[496] = 10'h05f;
        mem[497] = 10'h283;
        mem[498] = 10'h2e7;
        mem[499] = 10'h2f9;
        mem[500] = 10'h318;
        mem[501] = 10'h112;
        mem[502] = 10'h3d8;
        mem[503] = 10'h068;
        mem[504] = 10'h13b;
        mem[505] = 10'h10a;
        mem[506] = 10'h281;
        mem[507] = 10'h0d1;
        mem[508] = 10'h3be;
        mem[509] = 10'h118;
        mem[510] = 10'h15b;
        mem[511] = 10'h2f2;
        mem[512] = 10'h0bd;
        mem[513] = 10'h1d9;
        mem[514] = 10'h16e;
        mem[515] = 10'h13c;
        mem[516] = 10'h34b;
        mem[517] = 10'h005;
        mem[518] = 10'h334;
        mem[519] = 10'h173;
        mem[520] = 10'h084;
        mem[521] = 10'h030;
        mem[522] = 10'h311;
        mem[523] = 10'h0d5;
        mem[524] = 10'h393;
        mem[525] = 10'h01a;
        mem[526] = 10'h36f;
        mem[527] = 10'h230;
        mem[528] = 10'h174;
        mem[529] = 10'h11e;
        mem[530] = 10'h02a;
        mem[531] = 10'h27e;
        mem[532] = 10'h363;
        mem[533] = 10'h39f;
        mem[534] = 10'h116;
        mem[535] = 10'h287;
        mem[536] = 10'h1bf;
        mem[537] = 10'h3ed;
        mem[538] = 10'h0d6;
        mem[539] = 10'h2bf;
        mem[540] = 10'h2ba;
        mem[541] = 10'h087;
        mem[542] = 10'h12e;
        mem[543] = 10'h04e;
        mem[544] = 10'h154;
        mem[545] = 10'h01f;
        mem[546] = 10'h224;
        mem[547] = 10'h358;
        mem[548] = 10'h3ef;
        mem[549] = 10'h0d8;
        mem[550] = 10'h1e7;
        mem[551] = 10'h0b2;
        mem[552] = 10'h0d9;
        mem[553] = 10'h2e4;
        mem[554] = 10'h1f4;
        mem[555] = 10'h38b;
        mem[556] = 10'h2e5;
        mem[557] = 10'h040;
        mem[558] = 10'h08e;
        mem[559] = 10'h325;
        mem[560] = 10'h2a7;
        mem[561] = 10'h38c;
        mem[562] = 10'h24f;
        mem[563] = 10'h143;
        mem[564] = 10'h12a;
        mem[565] = 10'h34a;
        mem[566] = 10'h02b;
        mem[567] = 10'h357;
        mem[568] = 10'h2ac;
        mem[569] = 10'h2d7;
        mem[570] = 10'h09f;
        mem[571] = 10'h35d;
        mem[572] = 10'h186;
        mem[573] = 10'h1d1;
        mem[574] = 10'h1e9;
        mem[575] = 10'h04b;
        mem[576] = 10'h126;
        mem[577] = 10'h332;
        mem[578] = 10'h2ef;
        mem[579] = 10'h1c3;
        mem[580] = 10'h034;
        mem[581] = 10'h35f;
        mem[582] = 10'h1d0;
        mem[583] = 10'h324;
        mem[584] = 10'h10f;
        mem[585] = 10'h298;
        mem[586] = 10'h0e1;
        mem[587] = 10'h2c6;
        mem[588] = 10'h222;
        mem[589] = 10'h3c1;
        mem[590] = 10'h23f;
        mem[591] = 10'h004;
        mem[592] = 10'h169;
        mem[593] = 10'h1f2;
        mem[594] = 10'h2ec;
        mem[595] = 10'h36d;
        mem[596] = 10'h18a;
        mem[597] = 10'h0ba;
        mem[598] = 10'h221;
        mem[599] = 10'h33d;
        mem[600] = 10'h39a;
        mem[601] = 10'h2c9;
        mem[602] = 10'h0aa;
        mem[603] = 10'h1a9;
        mem[604] = 10'h30a;
        mem[605] = 10'h083;
        mem[606] = 10'h2c5;
        mem[607] = 10'h3db;
        mem[608] = 10'h196;
        mem[609] = 10'h203;
        mem[610] = 10'h341;
        mem[611] = 10'h30e;
        mem[612] = 10'h389;
        mem[613] = 10'h2b5;
        mem[614] = 10'h00a;
        mem[615] = 10'h082;
        mem[616] = 10'h014;
        mem[617] = 10'h02f;
        mem[618] = 10'h3da;
        mem[619] = 10'h0f5;
        mem[620] = 10'h295;
        mem[621] = 10'h241;
        mem[622] = 10'h06d;
        mem[623] = 10'h269;
        mem[624] = 10'h264;
        mem[625] = 10'h05d;
        mem[626] = 10'h3a5;
        mem[627] = 10'h1b5;
        mem[628] = 10'h3e6;
        mem[629] = 10'h2ea;
        mem[630] = 10'h0b3;
        mem[631] = 10'h1f9;
        mem[632] = 10'h00e;
        mem[633] = 10'h170;
        mem[634] = 10'h1de;
        mem[635] = 10'h3ff;
        mem[636] = 10'h0b7;
        mem[637] = 10'h275;
        mem[638] = 10'h320;
        mem[639] = 10'h0e5;
        mem[640] = 10'h0e2;
        mem[641] = 10'h243;
        mem[642] = 10'h16b;
        mem[643] = 10'h33b;
        mem[644] = 10'h048;
        mem[645] = 10'h1d8;
        mem[646] = 10'h252;
        mem[647] = 10'h3b4;
        mem[648] = 10'h3f1;
        mem[649] = 10'h0fc;
        mem[650] = 10'h2c3;
        mem[651] = 10'h30f;
        mem[652] = 10'h28e;
        mem[653] = 10'h316;
        mem[654] = 10'h0eb;
        mem[655] = 10'h3e0;
        mem[656] = 10'h360;
        mem[657] = 10'h0cc;
        mem[658] = 10'h070;
        mem[659] = 10'h36b;
        mem[660] = 10'h25d;
        mem[661] = 10'h2b0;
        mem[662] = 10'h103;
        mem[663] = 10'h097;
        mem[664] = 10'h3f9;
        mem[665] = 10'h303;
        mem[666] = 10'h14d;
        mem[667] = 10'h130;
        mem[668] = 10'h3f5;
        mem[669] = 10'h10e;
        mem[670] = 10'h188;
        mem[671] = 10'h218;
        mem[672] = 10'h3ea;
        mem[673] = 10'h145;
        mem[674] = 10'h3e9;
        mem[675] = 10'h255;
        mem[676] = 10'h3a2;
        mem[677] = 10'h056;
        mem[678] = 10'h1fc;
        mem[679] = 10'h2f6;
        mem[680] = 10'h0e3;
        mem[681] = 10'h19d;
        mem[682] = 10'h326;
        mem[683] = 10'h25c;
        mem[684] = 10'h047;
        mem[685] = 10'h197;
        mem[686] = 10'h3b9;
        mem[687] = 10'h210;
        mem[688] = 10'h1d4;
        mem[689] = 10'h261;
        mem[690] = 10'h2b2;
        mem[691] = 10'h3ba;
        mem[692] = 10'h100;
        mem[693] = 10'h3c2;
        mem[694] = 10'h3ca;
        mem[695] = 10'h0f8;
        mem[696] = 10'h277;
        mem[697] = 10'h028;
        mem[698] = 10'h0af;
        mem[699] = 10'h10d;
        mem[700] = 10'h2d8;
        mem[701] = 10'h273;
        mem[702] = 10'h101;
        mem[703] = 10'h3f2;
        mem[704] = 10'h15f;
        mem[705] = 10'h05c;
        mem[706] = 10'h0be;
        mem[707] = 10'h2f3;
        mem[708] = 10'h0a8;
        mem[709] = 10'h136;
        mem[710] = 10'h0e0;
        mem[711] = 10'h01b;
        mem[712] = 10'h373;
        mem[713] = 10'h3cf;
        mem[714] = 10'h370;
        mem[715] = 10'h148;
        mem[716] = 10'h03d;
        mem[717] = 10'h138;
        mem[718] = 10'h362;
        mem[719] = 10'h2e6;
        mem[720] = 10'h07f;
        mem[721] = 10'h366;
        mem[722] = 10'h32c;
        mem[723] = 10'h190;
        mem[724] = 10'h346;
        mem[725] = 10'h0ef;
        mem[726] = 10'h0ad;
        mem[727] = 10'h33a;
        mem[728] = 10'h30d;
        mem[729] = 10'h171;
        mem[730] = 10'h3c0;
        mem[731] = 10'h17c;
        mem[732] = 10'h280;
        mem[733] = 10'h009;
        mem[734] = 10'h2d9;
        mem[735] = 10'h023;
        mem[736] = 10'h092;
        mem[737] = 10'h2ce;
        mem[738] = 10'h3bf;
        mem[739] = 10'h1d7;
        mem[740] = 10'h146;
        mem[741] = 10'h155;
        mem[742] = 10'h20d;
        mem[743] = 10'h160;
        mem[744] = 10'h168;
        mem[745] = 10'h3d1;
        mem[746] = 10'h172;
        mem[747] = 10'h1a6;
        mem[748] = 10'h01e;
        mem[749] = 10'h3a8;
        mem[750] = 10'h37a;
        mem[751] = 10'h2d3;
        mem[752] = 10'h240;
        mem[753] = 10'h03a;
        mem[754] = 10'h259;
        mem[755] = 10'h06a;
        mem[756] = 10'h2fa;
        mem[757] = 10'h0b8;
        mem[758] = 10'h0fe;
        mem[759] = 10'h361;
        mem[760] = 10'h3ee;
        mem[761] = 10'h249;
        mem[762] = 10'h00f;
        mem[763] = 10'h20a;
        mem[764] = 10'h0a5;
        mem[765] = 10'h010;
        mem[766] = 10'h200;
        mem[767] = 10'h2f1;
        mem[768] = 10'h0bf;
        mem[769] = 10'h1ec;
        mem[770] = 10'h06b;
        mem[771] = 10'h2cd;
        mem[772] = 10'h2da;
        mem[773] = 10'h1a7;
        mem[774] = 10'h365;
        mem[775] = 10'h314;
        mem[776] = 10'h3ad;
        mem[777] = 10'h1b3;
        mem[778] = 10'h0f0;
        mem[779] = 10'h1ca;
        mem[780] = 10'h25e;
        mem[781] = 10'h043;
        mem[782] = 10'h214;
        mem[783] = 10'h04c;
        mem[784] = 10'h2d5;
        mem[785] = 10'h14a;
        mem[786] = 10'h2ff;
        mem[787] = 10'h0d3;
        mem[788] = 10'h2a6;
        mem[789] = 10'h179;
        mem[790] = 10'h0ec;
        mem[791] = 10'h150;
        mem[792] = 10'h181;
        mem[793] = 10'h175;
        mem[794] = 10'h3a1;
        mem[795] = 10'h1bb;
        mem[796] = 10'h253;
        mem[797] = 10'h356;
        mem[798] = 10'h3dd;
        mem[799] = 10'h2cc;
        mem[800] = 10'h38a;
        mem[801] = 10'h396;
        mem[802] = 10'h2dc;
        mem[803] = 10'h122;
        mem[804] = 10'h3f6;
        mem[805] = 10'h23c;
        mem[806] = 10'h18d;
        mem[807] = 10'h248;
        mem[808] = 10'h382;
        mem[809] = 10'h2ca;
        mem[810] = 10'h239;
        mem[811] = 10'h1a0;
        mem[812] = 10'h2e9;
        mem[813] = 10'h15d;
        mem[814] = 10'h3dc;
        mem[815] = 10'h099;
        mem[816] = 10'h026;
        mem[817] = 10'h05a;
        mem[818] = 10'h098;
        mem[819] = 10'h2d0;
        mem[820] = 10'h247;
        mem[821] = 10'h37f;
        mem[822] = 10'h25f;
        mem[823] = 10'h104;
        mem[824] = 10'h1f6;
        mem[825] = 10'h2bd;
        mem[826] = 10'h194;
        mem[827] = 10'h1aa;
        mem[828] = 10'h198;
        mem[829] = 10'h165;
        mem[830] = 10'h270;
        mem[831] = 10'h0cb;
        mem[832] = 10'h177;
        mem[833] = 10'h2a5;
        mem[834] = 10'h2bb;
        mem[835] = 10'h015;
        mem[836] = 10'h371;
        mem[837] = 10'h2c4;
        mem[838] = 10'h132;
        mem[839] = 10'h323;
        mem[840] = 10'h385;
        mem[841] = 10'h16f;
        mem[842] = 10'h153;
        mem[843] = 10'h3ae;
        mem[844] = 10'h3d4;
        mem[845] = 10'h1f5;
        mem[846] = 10'h0c0;
        mem[847] = 10'h206;
        mem[848] = 10'h17a;
        mem[849] = 10'h23d;
        mem[850] = 10'h3e7;
        mem[851] = 10'h00d;
        mem[852] = 10'h069;
        mem[853] = 10'h322;
        mem[854] = 10'h3eb;
        mem[855] = 10'h1a4;
        mem[856] = 10'h3a0;
        mem[857] = 10'h23a;
        mem[858] = 10'h17b;
        mem[859] = 10'h096;
        mem[860] = 10'h18e;
        mem[861] = 10'h07d;
        mem[862] = 10'h09e;
        mem[863] = 10'h0bc;
        mem[864] = 10'h304;
        mem[865] = 10'h21d;
        mem[866] = 10'h135;
        mem[867] = 10'h267;
        mem[868] = 10'h192;
        mem[869] = 10'h066;
        mem[870] = 10'h384;
        mem[871] = 10'h12f;
        mem[872] = 10'h1ba;
        mem[873] = 10'h232;
        mem[874] = 10'h0a7;
        mem[875] = 10'h34d;
        mem[876] = 10'h288;
        mem[877] = 10'h163;
        mem[878] = 10'h0c1;
        mem[879] = 10'h2ed;
        mem[880] = 10'h20c;
        mem[881] = 10'h381;
        mem[882] = 10'h091;
        mem[883] = 10'h3f3;
        mem[884] = 10'h03c;
        mem[885] = 10'h02c;
        mem[886] = 10'h282;
        mem[887] = 10'h19a;
        mem[888] = 10'h185;
        mem[889] = 10'h211;
        mem[890] = 10'h351;
        mem[891] = 10'h178;
        mem[892] = 10'h21b;
        mem[893] = 10'h07e;
        mem[894] = 10'h37b;
        mem[895] = 10'h2f7;
        mem[896] = 10'h226;
        mem[897] = 10'h22c;
        mem[898] = 10'h1e1;
        mem[899] = 10'h0f3;
        mem[900] = 10'h128;
        mem[901] = 10'h27b;
        mem[902] = 10'h1d3;
        mem[903] = 10'h1bd;
        mem[904] = 10'h0fa;
        mem[905] = 10'h1c7;
        mem[906] = 10'h2a1;
        mem[907] = 10'h3c8;
        mem[908] = 10'h31c;
        mem[909] = 10'h31d;
        mem[910] = 10'h38d;
        mem[911] = 10'h2d4;
        mem[912] = 10'h32b;
        mem[913] = 10'h3e2;
        mem[914] = 10'h265;
        mem[915] = 10'h354;
        mem[916] = 10'h1d6;
        mem[917] = 10'h193;
        mem[918] = 10'h011;
        mem[919] = 10'h11a;
        mem[920] = 10'h233;
        mem[921] = 10'h23b;
        mem[922] = 10'h3f7;
        mem[923] = 10'h392;
        mem[924] = 10'h1ed;
        mem[925] = 10'h327;
        mem[926] = 10'h367;
        mem[927] = 10'h144;
        mem[928] = 10'h33c;
        mem[929] = 10'h2a3;
        mem[930] = 10'h319;
        mem[931] = 10'h1fa;
        mem[932] = 10'h300;
        mem[933] = 10'h374;
        mem[934] = 10'h3bc;
        mem[935] = 10'h021;
        mem[936] = 10'h183;
        mem[937] = 10'h397;
        mem[938] = 10'h04d;
        mem[939] = 10'h09d;
        mem[940] = 10'h036;
        mem[941] = 10'h29e;
        mem[942] = 10'h29d;
        mem[943] = 10'h250;
        mem[944] = 10'h1c2;
        mem[945] = 10'h2aa;
        mem[946] = 10'h290;
        mem[947] = 10'h127;
        mem[948] = 10'h289;
        mem[949] = 10'h032;
        mem[950] = 10'h378;
        mem[951] = 10'h184;
        mem[952] = 10'h237;
        mem[953] = 10'h2bc;
        mem[954] = 10'h22d;
        mem[955] = 10'h0a1;
        mem[956] = 10'h139;
        mem[957] = 10'h0f2;
        mem[958] = 10'h3ce;
        mem[959] = 10'h1f8;
        mem[960] = 10'h2dd;
        mem[961] = 10'h3d3;
        mem[962] = 10'h3d6;
        mem[963] = 10'h031;
        mem[964] = 10'h0dc;
        mem[965] = 10'h3bd;
        mem[966] = 10'h1e5;
        mem[967] = 10'h28a;
        mem[968] = 10'h3b1;
        mem[969] = 10'h012;
        mem[970] = 10'h1cb;
        mem[971] = 10'h3c4;
        mem[972] = 10'h16d;
        mem[973] = 10'h01c;
        mem[974] = 10'h345;
        mem[975] = 10'h234;
        mem[976] = 10'h13e;
        mem[977] = 10'h018;
        mem[978] = 10'h2ae;
        mem[979] = 10'h375;
        mem[980] = 10'h086;
        mem[981] = 10'h003;
        mem[982] = 10'h0b4;
        mem[983] = 10'h29f;
        mem[984] = 10'h20e;
        mem[985] = 10'h074;
        mem[986] = 10'h379;
        mem[987] = 10'h07b;
        mem[988] = 10'h29a;
        mem[989] = 10'h26d;
        mem[990] = 10'h235;
        mem[991] = 10'h399;
        mem[992] = 10'h0bb;
        mem[993] = 10'h1fe;
        mem[994] = 10'h17e;
        mem[995] = 10'h27a;
        mem[996] = 10'h113;
        mem[997] = 10'h062;
        mem[998] = 10'h1ae;
        mem[999] = 10'h025;
        mem[1000] = 10'h24b;
        mem[1001] = 10'h072;
        mem[1002] = 10'h246;
        mem[1003] = 10'h0b9;
        mem[1004] = 10'h328;
        mem[1005] = 10'h228;
        mem[1006] = 10'h079;
        mem[1007] = 10'h020;
        mem[1008] = 10'h2d6;
        mem[1009] = 10'h220;
        mem[1010] = 10'h3a3;
        mem[1011] = 10'h219;
        mem[1012] = 10'h35e;
        mem[1013] = 10'h376;
        mem[1014] = 10'h15c;
        mem[1015] = 10'h076;
        mem[1016] = 10'h14e;
        mem[1017] = 10'h027;
        mem[1018] = 10'h065;
        mem[1019] = 10'h3af;
        mem[1020] = 10'h1ff;
        mem[1021] = 10'h04f;
        mem[1022] = 10'h073;
        mem[1023] = 10'h1dc;
    end
endmodule

module odo_sbox_large2(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h161;
        mem[1] = 10'h270;
        mem[2] = 10'h38d;
        mem[3] = 10'h398;
        mem[4] = 10'h023;
        mem[5] = 10'h2a8;
        mem[6] = 10'h116;
        mem[7] = 10'h303;
        mem[8] = 10'h24a;
        mem[9] = 10'h0d3;
        mem[10] = 10'h18d;
        mem[11] = 10'h190;
        mem[12] = 10'h284;
        mem[13] = 10'h372;
        mem[14] = 10'h1de;
        mem[15] = 10'h3f7;
        mem[16] = 10'h21d;
        mem[17] = 10'h0bb;
        mem[18] = 10'h3fb;
        mem[19] = 10'h096;
        mem[20] = 10'h02c;
        mem[21] = 10'h130;
        mem[22] = 10'h1eb;
        mem[23] = 10'h339;
        mem[24] = 10'h391;
        mem[25] = 10'h2a6;
        mem[26] = 10'h082;
        mem[27] = 10'h3c7;
        mem[28] = 10'h315;
        mem[29] = 10'h183;
        mem[30] = 10'h143;
        mem[31] = 10'h0de;
        mem[32] = 10'h235;
        mem[33] = 10'h181;
        mem[34] = 10'h04d;
        mem[35] = 10'h32e;
        mem[36] = 10'h3f5;
        mem[37] = 10'h0dd;
        mem[38] = 10'h122;
        mem[39] = 10'h008;
        mem[40] = 10'h227;
        mem[41] = 10'h215;
        mem[42] = 10'h334;
        mem[43] = 10'h17c;
        mem[44] = 10'h0f6;
        mem[45] = 10'h050;
        mem[46] = 10'h13f;
        mem[47] = 10'h100;
        mem[48] = 10'h3fc;
        mem[49] = 10'h355;
        mem[50] = 10'h049;
        mem[51] = 10'h152;
        mem[52] = 10'h063;
        mem[53] = 10'h3d5;
        mem[54] = 10'h3b5;
        mem[55] = 10'h21f;
        mem[56] = 10'h24e;
        mem[57] = 10'h35b;
        mem[58] = 10'h185;
        mem[59] = 10'h094;
        mem[60] = 10'h1fa;
        mem[61] = 10'h1c8;
        mem[62] = 10'h2d6;
        mem[63] = 10'h12c;
        mem[64] = 10'h2f4;
        mem[65] = 10'h1f0;
        mem[66] = 10'h0c1;
        mem[67] = 10'h14f;
        mem[68] = 10'h218;
        mem[69] = 10'h1dd;
        mem[70] = 10'h00d;
        mem[71] = 10'h163;
        mem[72] = 10'h097;
        mem[73] = 10'h2ca;
        mem[74] = 10'h20e;
        mem[75] = 10'h057;
        mem[76] = 10'h39e;
        mem[77] = 10'h3fd;
        mem[78] = 10'h306;
        mem[79] = 10'h261;
        mem[80] = 10'h3ec;
        mem[81] = 10'h0c2;
        mem[82] = 10'h151;
        mem[83] = 10'h38c;
        mem[84] = 10'h295;
        mem[85] = 10'h3f8;
        mem[86] = 10'h3c6;
        mem[87] = 10'h2af;
        mem[88] = 10'h3ed;
        mem[89] = 10'h3af;
        mem[90] = 10'h20d;
        mem[91] = 10'h17a;
        mem[92] = 10'h093;
        mem[93] = 10'h3e4;
        mem[94] = 10'h393;
        mem[95] = 10'h3d9;
        mem[96] = 10'h18b;
        mem[97] = 10'h3a6;
        mem[98] = 10'h188;
        mem[99] = 10'h006;
        mem[100] = 10'h0a9;
        mem[101] = 10'h060;
        mem[102] = 10'h073;
        mem[103] = 10'h06a;
        mem[104] = 10'h01b;
        mem[105] = 10'h327;
        mem[106] = 10'h254;
        mem[107] = 10'h026;
        mem[108] = 10'h338;
        mem[109] = 10'h2ae;
        mem[110] = 10'h27b;
        mem[111] = 10'h102;
        mem[112] = 10'h0f0;
        mem[113] = 10'h167;
        mem[114] = 10'h2bb;
        mem[115] = 10'h089;
        mem[116] = 10'h353;
        mem[117] = 10'h029;
        mem[118] = 10'h366;
        mem[119] = 10'h27c;
        mem[120] = 10'h12e;
        mem[121] = 10'h3e7;
        mem[122] = 10'h02e;
        mem[123] = 10'h032;
        mem[124] = 10'h1a9;
        mem[125] = 10'h1a4;
        mem[126] = 10'h341;
        mem[127] = 10'h1ba;
        mem[128] = 10'h267;
        mem[129] = 10'h007;
        mem[130] = 10'h12a;
        mem[131] = 10'h0fa;
        mem[132] = 10'h24b;
        mem[133] = 10'h31e;
        mem[134] = 10'h3d7;
        mem[135] = 10'h140;
        mem[136] = 10'h076;
        mem[137] = 10'h0b9;
        mem[138] = 10'h1ae;
        mem[139] = 10'h1e2;
        mem[140] = 10'h0af;
        mem[141] = 10'h110;
        mem[142] = 10'h0e3;
        mem[143] = 10'h314;
        mem[144] = 10'h3e5;
        mem[145] = 10'h368;
        mem[146] = 10'h3a1;
        mem[147] = 10'h216;
        mem[148] = 10'h10a;
        mem[149] = 10'h0d6;
        mem[150] = 10'h179;
        mem[151] = 10'h149;
        mem[152] = 10'h15c;
        mem[153] = 10'h223;
        mem[154] = 10'h15d;
        mem[155] = 10'h27e;
        mem[156] = 10'h2f9;
        mem[157] = 10'h04c;
        mem[158] = 10'h3bb;
        mem[159] = 10'h287;
        mem[160] = 10'h0c8;
        mem[161] = 10'h275;
        mem[162] = 10'h241;
        mem[163] = 10'h268;
        mem[164] = 10'h3dc;
        mem[165] = 10'h033;
        mem[166] = 10'h36d;
        mem[167] = 10'h376;
        mem[168] = 10'h321;
        mem[169] = 10'h0bf;
        mem[170] = 10'h2f2;
        mem[171] = 10'h020;
        mem[172] = 10'h2f0;
        mem[173] = 10'h194;
        mem[174] = 10'h028;
        mem[175] = 10'h207;
        mem[176] = 10'h2df;
        mem[177] = 10'h2d3;
        mem[178] = 10'h1f1;
        mem[179] = 10'h0fc;
        mem[180] = 10'h329;
        mem[181] = 10'h1ce;
        mem[182] = 10'h040;
        mem[183] = 10'h072;
        mem[184] = 10'h210;
        mem[185] = 10'h09a;
        mem[186] = 10'h3bf;
        mem[187] = 10'h08c;
        mem[188] = 10'h05c;
        mem[189] = 10'h3b9;
        mem[190] = 10'h20a;
        mem[191] = 10'h024;
        mem[192] = 10'h004;
        mem[193] = 10'h035;
        mem[194] = 10'h2cb;
        mem[195] = 10'h3e6;
        mem[196] = 10'h390;
        mem[197] = 10'h3f2;
        mem[198] = 10'h3b3;
        mem[199] = 10'h1fc;
        mem[200] = 10'h2e9;
        mem[201] = 10'h30a;
        mem[202] = 10'h277;
        mem[203] = 10'h37e;
        mem[204] = 10'h0f8;
        mem[205] = 10'h1db;
        mem[206] = 10'h155;
        mem[207] = 10'h3a2;
        mem[208] = 10'h1d8;
        mem[209] = 10'h1fd;
        mem[210] = 10'h126;
        mem[211] = 10'h3a4;
        mem[212] = 10'h0c9;
        mem[213] = 10'h153;
        mem[214] = 10'h285;
        mem[215] = 10'h087;
        mem[216] = 10'h2c0;
        mem[217] = 10'h00a;
        mem[218] = 10'h0a8;
        mem[219] = 10'h2c5;
        mem[220] = 10'h067;
        mem[221] = 10'h186;
        mem[222] = 10'h2b8;
        mem[223] = 10'h247;
        mem[224] = 10'h00c;
        mem[225] = 10'h15b;
        mem[226] = 10'h3eb;
        mem[227] = 10'h20f;
        mem[228] = 10'h0a0;
        mem[229] = 10'h0e2;
        mem[230] = 10'h2ec;
        mem[231] = 10'h313;
        mem[232] = 10'h2a0;
        mem[233] = 10'h225;
        mem[234] = 10'h290;
        mem[235] = 10'h1e6;
        mem[236] = 10'h123;
        mem[237] = 10'h3bc;
        mem[238] = 10'h16a;
        mem[239] = 10'h37a;
        mem[240] = 10'h219;
        mem[241] = 10'h28a;
        mem[242] = 10'h3f1;
        mem[243] = 10'h2a7;
        mem[244] = 10'h1b8;
        mem[245] = 10'h03b;
        mem[246] = 10'h33d;
        mem[247] = 10'h22b;
        mem[248] = 10'h168;
        mem[249] = 10'h17f;
        mem[250] = 10'h156;
        mem[251] = 10'h1da;
        mem[252] = 10'h03f;
        mem[253] = 10'h07c;
        mem[254] = 10'h26d;
        mem[255] = 10'h027;
        mem[256] = 10'h0dc;
        mem[257] = 10'h174;
        mem[258] = 10'h068;
        mem[259] = 10'h0b1;
        mem[260] = 10'h132;
        mem[261] = 10'h146;
        mem[262] = 10'h3c9;
        mem[263] = 10'h02d;
        mem[264] = 10'h2de;
        mem[265] = 10'h1b6;
        mem[266] = 10'h1b0;
        mem[267] = 10'h1cc;
        mem[268] = 10'h2fe;
        mem[269] = 10'h1fb;
        mem[270] = 10'h134;
        mem[271] = 10'h1d3;
        mem[272] = 10'h090;
        mem[273] = 10'h042;
        mem[274] = 10'h159;
        mem[275] = 10'h09c;
        mem[276] = 10'h1d7;
        mem[277] = 10'h30b;
        mem[278] = 10'h32d;
        mem[279] = 10'h08b;
        mem[280] = 10'h2d9;
        mem[281] = 10'h294;
        mem[282] = 10'h0c5;
        mem[283] = 10'h0d9;
        mem[284] = 10'h10b;
        mem[285] = 10'h0d0;
        mem[286] = 10'h2b2;
        mem[287] = 10'h045;
        mem[288] = 10'h25b;
        mem[289] = 10'h15f;
        mem[290] = 10'h091;
        mem[291] = 10'h25f;
        mem[292] = 10'h09b;
        mem[293] = 10'h3cc;
        mem[294] = 10'h133;
        mem[295] = 10'h382;
        mem[296] = 10'h2f6;
        mem[297] = 10'h3db;
        mem[298] = 10'h205;
        mem[299] = 10'h069;
        mem[300] = 10'h021;
        mem[301] = 10'h01a;
        mem[302] = 10'h065;
        mem[303] = 10'h0f4;
        mem[304] = 10'h0f9;
        mem[305] = 10'h0be;
        mem[306] = 10'h14a;
        mem[307] = 10'h375;
        mem[308] = 10'h242;
        mem[309] = 10'h39d;
        mem[310] = 10'h1c1;
        mem[311] = 10'h240;
        mem[312] = 10'h18c;
        mem[313] = 10'h080;
        mem[314] = 10'h26a;
        mem[315] = 10'h1ee;
        mem[316] = 10'h06c;
        mem[317] = 10'h05d;
        mem[318] = 10'h2ea;
        mem[319] = 10'h09e;
        mem[320] = 10'h374;
        mem[321] = 10'h113;
        mem[322] = 10'h0eb;
        mem[323] = 10'h148;
        mem[324] = 10'h1c0;
        mem[325] = 10'h0d1;
        mem[326] = 10'h27f;
        mem[327] = 10'h32a;
        mem[328] = 10'h3fe;
        mem[329] = 10'h1cd;
        mem[330] = 10'h002;
        mem[331] = 10'h139;
        mem[332] = 10'h05a;
        mem[333] = 10'h1cb;
        mem[334] = 10'h3ef;
        mem[335] = 10'h1f7;
        mem[336] = 10'h070;
        mem[337] = 10'h3ba;
        mem[338] = 10'h119;
        mem[339] = 10'h274;
        mem[340] = 10'h349;
        mem[341] = 10'h3c2;
        mem[342] = 10'h3e1;
        mem[343] = 10'h3de;
        mem[344] = 10'h2da;
        mem[345] = 10'h0e9;
        mem[346] = 10'h38b;
        mem[347] = 10'h005;
        mem[348] = 10'h016;
        mem[349] = 10'h286;
        mem[350] = 10'h095;
        mem[351] = 10'h150;
        mem[352] = 10'h02f;
        mem[353] = 10'h15e;
        mem[354] = 10'h138;
        mem[355] = 10'h1d1;
        mem[356] = 10'h012;
        mem[357] = 10'h3e8;
        mem[358] = 10'h3ee;
        mem[359] = 10'h288;
        mem[360] = 10'h1f3;
        mem[361] = 10'h202;
        mem[362] = 10'h32f;
        mem[363] = 10'h1ca;
        mem[364] = 10'h320;
        mem[365] = 10'h0ac;
        mem[366] = 10'h30c;
        mem[367] = 10'h030;
        mem[368] = 10'h3d3;
        mem[369] = 10'h196;
        mem[370] = 10'h3cd;
        mem[371] = 10'h0b0;
        mem[372] = 10'h37d;
        mem[373] = 10'h165;
        mem[374] = 10'h099;
        mem[375] = 10'h05b;
        mem[376] = 10'h3df;
        mem[377] = 10'h34e;
        mem[378] = 10'h377;
        mem[379] = 10'h332;
        mem[380] = 10'h2db;
        mem[381] = 10'h26e;
        mem[382] = 10'h0f7;
        mem[383] = 10'h192;
        mem[384] = 10'h3a7;
        mem[385] = 10'h0cd;
        mem[386] = 10'h1c7;
        mem[387] = 10'h02a;
        mem[388] = 10'h2e8;
        mem[389] = 10'h39f;
        mem[390] = 10'h182;
        mem[391] = 10'h3aa;
        mem[392] = 10'h370;
        mem[393] = 10'h191;
        mem[394] = 10'h2fd;
        mem[395] = 10'h025;
        mem[396] = 10'h0cb;
        mem[397] = 10'h2ad;
        mem[398] = 10'h09d;
        mem[399] = 10'h298;
        mem[400] = 10'h3c1;
        mem[401] = 10'h28f;
        mem[402] = 10'h3ad;
        mem[403] = 10'h0fe;
        mem[404] = 10'h098;
        mem[405] = 10'h324;
        mem[406] = 10'h23b;
        mem[407] = 10'h13e;
        mem[408] = 10'h251;
        mem[409] = 10'h104;
        mem[410] = 10'h2a9;
        mem[411] = 10'h0c3;
        mem[412] = 10'h2f7;
        mem[413] = 10'h24d;
        mem[414] = 10'h36b;
        mem[415] = 10'h3b0;
        mem[416] = 10'h2bd;
        mem[417] = 10'h27a;
        mem[418] = 10'h380;
        mem[419] = 10'h1e0;
        mem[420] = 10'h08f;
        mem[421] = 10'h3dd;
        mem[422] = 10'h171;
        mem[423] = 10'h041;
        mem[424] = 10'h11c;
        mem[425] = 10'h394;
        mem[426] = 10'h2d2;
        mem[427] = 10'h22f;
        mem[428] = 10'h33a;
        mem[429] = 10'h38e;
        mem[430] = 10'h2e3;
        mem[431] = 10'h058;
        mem[432] = 10'h363;
        mem[433] = 10'h056;
        mem[434] = 10'h1b4;
        mem[435] = 10'h112;
        mem[436] = 10'h193;
        mem[437] = 10'h301;
        mem[438] = 10'h21a;
        mem[439] = 10'h3b7;
        mem[440] = 10'h061;
        mem[441] = 10'h141;
        mem[442] = 10'h3ca;
        mem[443] = 10'h1bb;
        mem[444] = 10'h1c9;
        mem[445] = 10'h103;
        mem[446] = 10'h2be;
        mem[447] = 10'h051;
        mem[448] = 10'h083;
        mem[449] = 10'h1aa;
        mem[450] = 10'h231;
        mem[451] = 10'h378;
        mem[452] = 10'h160;
        mem[453] = 10'h20c;
        mem[454] = 10'h1c4;
        mem[455] = 10'h17e;
        mem[456] = 10'h316;
        mem[457] = 10'h2c8;
        mem[458] = 10'h044;
        mem[459] = 10'h1a6;
        mem[460] = 10'h35e;
        mem[461] = 10'h3d2;
        mem[462] = 10'h1a3;
        mem[463] = 10'h263;
        mem[464] = 10'h3f6;
        mem[465] = 10'h2cd;
        mem[466] = 10'h224;
        mem[467] = 10'h34b;
        mem[468] = 10'h1b9;
        mem[469] = 10'h213;
        mem[470] = 10'h1ad;
        mem[471] = 10'h2a5;
        mem[472] = 10'h272;
        mem[473] = 10'h1ff;
        mem[474] = 10'h198;
        mem[475] = 10'h1e1;
        mem[476] = 10'h1ac;
        mem[477] = 10'h23d;
        mem[478] = 10'h1af;
        mem[479] = 10'h2c3;
        mem[480] = 10'h212;
        mem[481] = 10'h266;
        mem[482] = 10'h289;
        mem[483] = 10'h175;
        mem[484] = 10'h107;
        mem[485] = 10'h10d;
        mem[486] = 10'h1d2;
        mem[487] = 10'h0e7;
        mem[488] = 10'h1e9;
        mem[489] = 10'h075;
        mem[490] = 10'h297;
        mem[491] = 10'h3f4;
        mem[492] = 10'h293;
        mem[493] = 10'h3e0;
        mem[494] = 10'h2b3;
        mem[495] = 10'h31c;
        mem[496] = 10'h03a;
        mem[497] = 10'h3c5;
        mem[498] = 10'h2d5;
        mem[499] = 10'h173;
        mem[500] = 10'h199;
        mem[501] = 10'h2c7;
        mem[502] = 10'h237;
        mem[503] = 10'h3f9;
        mem[504] = 10'h0cf;
        mem[505] = 10'h357;
        mem[506] = 10'h371;
        mem[507] = 10'h37f;
        mem[508] = 10'h124;
        mem[509] = 10'h311;
        mem[510] = 10'h200;
        mem[511] = 10'h3ae;
        mem[512] = 10'h2b6;
        mem[513] = 10'h06e;
        mem[514] = 10'h1ab;
        mem[515] = 10'h318;
        mem[516] = 10'h0b7;
        mem[517] = 10'h0e6;
        mem[518] = 10'h013;
        mem[519] = 10'h1c3;
        mem[520] = 10'h208;
        mem[521] = 10'h0d7;
        mem[522] = 10'h085;
        mem[523] = 10'h13b;
        mem[524] = 10'h1ef;
        mem[525] = 10'h31a;
        mem[526] = 10'h2f1;
        mem[527] = 10'h249;
        mem[528] = 10'h109;
        mem[529] = 10'h331;
        mem[530] = 10'h2b9;
        mem[531] = 10'h22e;
        mem[532] = 10'h2e7;
        mem[533] = 10'h2b1;
        mem[534] = 10'h11a;
        mem[535] = 10'h034;
        mem[536] = 10'h348;
        mem[537] = 10'h3f3;
        mem[538] = 10'h011;
        mem[539] = 10'h344;
        mem[540] = 10'h0ec;
        mem[541] = 10'h001;
        mem[542] = 10'h081;
        mem[543] = 10'h23e;
        mem[544] = 10'h358;
        mem[545] = 10'h2fa;
        mem[546] = 10'h246;
        mem[547] = 10'h3ff;
        mem[548] = 10'h121;
        mem[549] = 10'h229;
        mem[550] = 10'h0f2;
        mem[551] = 10'h3b1;
        mem[552] = 10'h2e1;
        mem[553] = 10'h2aa;
        mem[554] = 10'h259;
        mem[555] = 10'h236;
        mem[556] = 10'h01f;
        mem[557] = 10'h1c2;
        mem[558] = 10'h00b;
        mem[559] = 10'h12f;
        mem[560] = 10'h0c6;
        mem[561] = 10'h1d5;
        mem[562] = 10'h2d4;
        mem[563] = 10'h333;
        mem[564] = 10'h253;
        mem[565] = 10'h12b;
        mem[566] = 10'h19c;
        mem[567] = 10'h256;
        mem[568] = 10'h381;
        mem[569] = 10'h3c4;
        mem[570] = 10'h365;
        mem[571] = 10'h3bd;
        mem[572] = 10'h1b2;
        mem[573] = 10'h379;
        mem[574] = 10'h009;
        mem[575] = 10'h335;
        mem[576] = 10'h347;
        mem[577] = 10'h2b4;
        mem[578] = 10'h03d;
        mem[579] = 10'h074;
        mem[580] = 10'h33b;
        mem[581] = 10'h010;
        mem[582] = 10'h2a1;
        mem[583] = 10'h031;
        mem[584] = 10'h15a;
        mem[585] = 10'h117;
        mem[586] = 10'h05e;
        mem[587] = 10'h11b;
        mem[588] = 10'h3ac;
        mem[589] = 10'h24c;
        mem[590] = 10'h1ec;
        mem[591] = 10'h33f;
        mem[592] = 10'h022;
        mem[593] = 10'h038;
        mem[594] = 10'h257;
        mem[595] = 10'h36f;
        mem[596] = 10'h18e;
        mem[597] = 10'h2b5;
        mem[598] = 10'h0f3;
        mem[599] = 10'h234;
        mem[600] = 10'h3ab;
        mem[601] = 10'h1a2;
        mem[602] = 10'h048;
        mem[603] = 10'h19f;
        mem[604] = 10'h176;
        mem[605] = 10'h264;
        mem[606] = 10'h03c;
        mem[607] = 10'h05f;
        mem[608] = 10'h2d7;
        mem[609] = 10'h1b3;
        mem[610] = 10'h25d;
        mem[611] = 10'h36e;
        mem[612] = 10'h385;
        mem[613] = 10'h260;
        mem[614] = 10'h211;
        mem[615] = 10'h362;
        mem[616] = 10'h079;
        mem[617] = 10'h2dd;
        mem[618] = 10'h217;
        mem[619] = 10'h220;
        mem[620] = 10'h064;
        mem[621] = 10'h354;
        mem[622] = 10'h2d0;
        mem[623] = 10'h0e8;
        mem[624] = 10'h32c;
        mem[625] = 10'h0ab;
        mem[626] = 10'h399;
        mem[627] = 10'h1a5;
        mem[628] = 10'h145;
        mem[629] = 10'h312;
        mem[630] = 10'h30e;
        mem[631] = 10'h3e2;
        mem[632] = 10'h197;
        mem[633] = 10'h092;
        mem[634] = 10'h2a3;
        mem[635] = 10'h106;
        mem[636] = 10'h2ce;
        mem[637] = 10'h19b;
        mem[638] = 10'h0ef;
        mem[639] = 10'h1ed;
        mem[640] = 10'h300;
        mem[641] = 10'h396;
        mem[642] = 10'h0f5;
        mem[643] = 10'h39a;
        mem[644] = 10'h23c;
        mem[645] = 10'h0d4;
        mem[646] = 10'h3d6;
        mem[647] = 10'h28c;
        mem[648] = 10'h3c8;
        mem[649] = 10'h39b;
        mem[650] = 10'h2c2;
        mem[651] = 10'h397;
        mem[652] = 10'h23f;
        mem[653] = 10'h255;
        mem[654] = 10'h052;
        mem[655] = 10'h14d;
        mem[656] = 10'h0f1;
        mem[657] = 10'h17d;
        mem[658] = 10'h16f;
        mem[659] = 10'h204;
        mem[660] = 10'h2bc;
        mem[661] = 10'h28e;
        mem[662] = 10'h282;
        mem[663] = 10'h06b;
        mem[664] = 10'h39c;
        mem[665] = 10'h1f6;
        mem[666] = 10'h292;
        mem[667] = 10'h2c6;
        mem[668] = 10'h350;
        mem[669] = 10'h137;
        mem[670] = 10'h279;
        mem[671] = 10'h305;
        mem[672] = 10'h21c;
        mem[673] = 10'h1a8;
        mem[674] = 10'h373;
        mem[675] = 10'h164;
        mem[676] = 10'h326;
        mem[677] = 10'h184;
        mem[678] = 10'h11e;
        mem[679] = 10'h017;
        mem[680] = 10'h14e;
        mem[681] = 10'h0b4;
        mem[682] = 10'h0b2;
        mem[683] = 10'h2cf;
        mem[684] = 10'h265;
        mem[685] = 10'h248;
        mem[686] = 10'h16b;
        mem[687] = 10'h066;
        mem[688] = 10'h195;
        mem[689] = 10'h2ff;
        mem[690] = 10'h1ea;
        mem[691] = 10'h276;
        mem[692] = 10'h129;
        mem[693] = 10'h252;
        mem[694] = 10'h13a;
        mem[695] = 10'h0ff;
        mem[696] = 10'h340;
        mem[697] = 10'h22c;
        mem[698] = 10'h054;
        mem[699] = 10'h203;
        mem[700] = 10'h280;
        mem[701] = 10'h059;
        mem[702] = 10'h187;
        mem[703] = 10'h0d2;
        mem[704] = 10'h086;
        mem[705] = 10'h000;
        mem[706] = 10'h383;
        mem[707] = 10'h19e;
        mem[708] = 10'h34d;
        mem[709] = 10'h26b;
        mem[710] = 10'h23a;
        mem[711] = 10'h0c0;
        mem[712] = 10'h384;
        mem[713] = 10'h07a;
        mem[714] = 10'h1a1;
        mem[715] = 10'h262;
        mem[716] = 10'h2d8;
        mem[717] = 10'h09f;
        mem[718] = 10'h16e;
        mem[719] = 10'h1d6;
        mem[720] = 10'h1bf;
        mem[721] = 10'h0fb;
        mem[722] = 10'h3a0;
        mem[723] = 10'h07e;
        mem[724] = 10'h0bc;
        mem[725] = 10'h21e;
        mem[726] = 10'h1c6;
        mem[727] = 10'h2f5;
        mem[728] = 10'h108;
        mem[729] = 10'h2e5;
        mem[730] = 10'h01c;
        mem[731] = 10'h01e;
        mem[732] = 10'h302;
        mem[733] = 10'h307;
        mem[734] = 10'h367;
        mem[735] = 10'h2bf;
        mem[736] = 10'h11f;
        mem[737] = 10'h0db;
        mem[738] = 10'h3a9;
        mem[739] = 10'h243;
        mem[740] = 10'h319;
        mem[741] = 10'h046;
        mem[742] = 10'h18a;
        mem[743] = 10'h3b2;
        mem[744] = 10'h04b;
        mem[745] = 10'h162;
        mem[746] = 10'h13c;
        mem[747] = 10'h228;
        mem[748] = 10'h0ad;
        mem[749] = 10'h06d;
        mem[750] = 10'h291;
        mem[751] = 10'h127;
        mem[752] = 10'h2ac;
        mem[753] = 10'h22a;
        mem[754] = 10'h1dc;
        mem[755] = 10'h158;
        mem[756] = 10'h201;
        mem[757] = 10'h1f2;
        mem[758] = 10'h304;
        mem[759] = 10'h3b6;
        mem[760] = 10'h22d;
        mem[761] = 10'h078;
        mem[762] = 10'h24f;
        mem[763] = 10'h0b5;
        mem[764] = 10'h28d;
        mem[765] = 10'h2eb;
        mem[766] = 10'h2ab;
        mem[767] = 10'h1be;
        mem[768] = 10'h33c;
        mem[769] = 10'h35d;
        mem[770] = 10'h33e;
        mem[771] = 10'h08a;
        mem[772] = 10'h258;
        mem[773] = 10'h1f9;
        mem[774] = 10'h0d8;
        mem[775] = 10'h105;
        mem[776] = 10'h3ea;
        mem[777] = 10'h2ed;
        mem[778] = 10'h0ea;
        mem[779] = 10'h29e;
        mem[780] = 10'h392;
        mem[781] = 10'h0da;
        mem[782] = 10'h19a;
        mem[783] = 10'h1bc;
        mem[784] = 10'h34c;
        mem[785] = 10'h3a8;
        mem[786] = 10'h2a2;
        mem[787] = 10'h3f0;
        mem[788] = 10'h1a0;
        mem[789] = 10'h206;
        mem[790] = 10'h2b7;
        mem[791] = 10'h323;
        mem[792] = 10'h1c5;
        mem[793] = 10'h245;
        mem[794] = 10'h36a;
        mem[795] = 10'h271;
        mem[796] = 10'h0ae;
        mem[797] = 10'h115;
        mem[798] = 10'h0d5;
        mem[799] = 10'h0a5;
        mem[800] = 10'h351;
        mem[801] = 10'h2fc;
        mem[802] = 10'h07d;
        mem[803] = 10'h31d;
        mem[804] = 10'h07f;
        mem[805] = 10'h395;
        mem[806] = 10'h018;
        mem[807] = 10'h2e6;
        mem[808] = 10'h35a;
        mem[809] = 10'h16c;
        mem[810] = 10'h2ee;
        mem[811] = 10'h142;
        mem[812] = 10'h317;
        mem[813] = 10'h07b;
        mem[814] = 10'h1e4;
        mem[815] = 10'h120;
        mem[816] = 10'h0e1;
        mem[817] = 10'h0a4;
        mem[818] = 10'h3c3;
        mem[819] = 10'h387;
        mem[820] = 10'h1cf;
        mem[821] = 10'h2c4;
        mem[822] = 10'h088;
        mem[823] = 10'h221;
        mem[824] = 10'h361;
        mem[825] = 10'h25e;
        mem[826] = 10'h0a7;
        mem[827] = 10'h3ce;
        mem[828] = 10'h144;
        mem[829] = 10'h2b0;
        mem[830] = 10'h3e3;
        mem[831] = 10'h003;
        mem[832] = 10'h34f;
        mem[833] = 10'h273;
        mem[834] = 10'h322;
        mem[835] = 10'h345;
        mem[836] = 10'h3e9;
        mem[837] = 10'h31f;
        mem[838] = 10'h238;
        mem[839] = 10'h3d8;
        mem[840] = 10'h36c;
        mem[841] = 10'h29f;
        mem[842] = 10'h111;
        mem[843] = 10'h2e4;
        mem[844] = 10'h281;
        mem[845] = 10'h20b;
        mem[846] = 10'h0bd;
        mem[847] = 10'h0a6;
        mem[848] = 10'h17b;
        mem[849] = 10'h3d0;
        mem[850] = 10'h1d4;
        mem[851] = 10'h014;
        mem[852] = 10'h3fa;
        mem[853] = 10'h169;
        mem[854] = 10'h2c9;
        mem[855] = 10'h0e5;
        mem[856] = 10'h35c;
        mem[857] = 10'h3a3;
        mem[858] = 10'h250;
        mem[859] = 10'h2a4;
        mem[860] = 10'h16d;
        mem[861] = 10'h0ca;
        mem[862] = 10'h02b;
        mem[863] = 10'h178;
        mem[864] = 10'h336;
        mem[865] = 10'h154;
        mem[866] = 10'h369;
        mem[867] = 10'h077;
        mem[868] = 10'h0c4;
        mem[869] = 10'h1e7;
        mem[870] = 10'h3cb;
        mem[871] = 10'h26f;
        mem[872] = 10'h2e0;
        mem[873] = 10'h13d;
        mem[874] = 10'h360;
        mem[875] = 10'h364;
        mem[876] = 10'h1d0;
        mem[877] = 10'h2dc;
        mem[878] = 10'h2e2;
        mem[879] = 10'h0c7;
        mem[880] = 10'h0ed;
        mem[881] = 10'h14c;
        mem[882] = 10'h039;
        mem[883] = 10'h053;
        mem[884] = 10'h084;
        mem[885] = 10'h125;
        mem[886] = 10'h214;
        mem[887] = 10'h1f4;
        mem[888] = 10'h0a3;
        mem[889] = 10'h328;
        mem[890] = 10'h2f8;
        mem[891] = 10'h3d1;
        mem[892] = 10'h308;
        mem[893] = 10'h1df;
        mem[894] = 10'h18f;
        mem[895] = 10'h03e;
        mem[896] = 10'h359;
        mem[897] = 10'h147;
        mem[898] = 10'h29d;
        mem[899] = 10'h26c;
        mem[900] = 10'h10e;
        mem[901] = 10'h2ba;
        mem[902] = 10'h309;
        mem[903] = 10'h19d;
        mem[904] = 10'h08d;
        mem[905] = 10'h0aa;
        mem[906] = 10'h04e;
        mem[907] = 10'h29c;
        mem[908] = 10'h055;
        mem[909] = 10'h209;
        mem[910] = 10'h3da;
        mem[911] = 10'h10f;
        mem[912] = 10'h135;
        mem[913] = 10'h283;
        mem[914] = 10'h2d1;
        mem[915] = 10'h38f;
        mem[916] = 10'h047;
        mem[917] = 10'h036;
        mem[918] = 10'h346;
        mem[919] = 10'h1fe;
        mem[920] = 10'h0e4;
        mem[921] = 10'h10c;
        mem[922] = 10'h3c0;
        mem[923] = 10'h172;
        mem[924] = 10'h0b6;
        mem[925] = 10'h230;
        mem[926] = 10'h25c;
        mem[927] = 10'h189;
        mem[928] = 10'h3b4;
        mem[929] = 10'h32b;
        mem[930] = 10'h1f8;
        mem[931] = 10'h3b8;
        mem[932] = 10'h14b;
        mem[933] = 10'h25a;
        mem[934] = 10'h1f5;
        mem[935] = 10'h06f;
        mem[936] = 10'h310;
        mem[937] = 10'h389;
        mem[938] = 10'h37b;
        mem[939] = 10'h043;
        mem[940] = 10'h1e5;
        mem[941] = 10'h04f;
        mem[942] = 10'h2ef;
        mem[943] = 10'h1e8;
        mem[944] = 10'h28b;
        mem[945] = 10'h30d;
        mem[946] = 10'h386;
        mem[947] = 10'h1b5;
        mem[948] = 10'h114;
        mem[949] = 10'h296;
        mem[950] = 10'h131;
        mem[951] = 10'h342;
        mem[952] = 10'h2cc;
        mem[953] = 10'h101;
        mem[954] = 10'h0b3;
        mem[955] = 10'h29b;
        mem[956] = 10'h222;
        mem[957] = 10'h01d;
        mem[958] = 10'h0e0;
        mem[959] = 10'h325;
        mem[960] = 10'h3a5;
        mem[961] = 10'h0b8;
        mem[962] = 10'h180;
        mem[963] = 10'h00e;
        mem[964] = 10'h11d;
        mem[965] = 10'h29a;
        mem[966] = 10'h0ee;
        mem[967] = 10'h00f;
        mem[968] = 10'h239;
        mem[969] = 10'h0cc;
        mem[970] = 10'h35f;
        mem[971] = 10'h37c;
        mem[972] = 10'h330;
        mem[973] = 10'h12d;
        mem[974] = 10'h1a7;
        mem[975] = 10'h177;
        mem[976] = 10'h38a;
        mem[977] = 10'h31b;
        mem[978] = 10'h062;
        mem[979] = 10'h21b;
        mem[980] = 10'h2c1;
        mem[981] = 10'h128;
        mem[982] = 10'h226;
        mem[983] = 10'h170;
        mem[984] = 10'h3be;
        mem[985] = 10'h1bd;
        mem[986] = 10'h2fb;
        mem[987] = 10'h1b7;
        mem[988] = 10'h2f3;
        mem[989] = 10'h34a;
        mem[990] = 10'h071;
        mem[991] = 10'h019;
        mem[992] = 10'h0df;
        mem[993] = 10'h1d9;
        mem[994] = 10'h27d;
        mem[995] = 10'h1b1;
        mem[996] = 10'h037;
        mem[997] = 10'h388;
        mem[998] = 10'h157;
        mem[999] = 10'h04a;
        mem[1000] = 10'h136;
        mem[1001] = 10'h278;
        mem[1002] = 10'h352;
        mem[1003] = 10'h166;
        mem[1004] = 10'h30f;
        mem[1005] = 10'h08e;
        mem[1006] = 10'h232;
        mem[1007] = 10'h3d4;
        mem[1008] = 10'h0a2;
        mem[1009] = 10'h0a1;
        mem[1010] = 10'h233;
        mem[1011] = 10'h0ba;
        mem[1012] = 10'h343;
        mem[1013] = 10'h1e3;
        mem[1014] = 10'h299;
        mem[1015] = 10'h3cf;
        mem[1016] = 10'h269;
        mem[1017] = 10'h015;
        mem[1018] = 10'h0ce;
        mem[1019] = 10'h337;
        mem[1020] = 10'h244;
        mem[1021] = 10'h356;
        mem[1022] = 10'h0fd;
        mem[1023] = 10'h118;
    end
endmodule

module odo_sbox_large3(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h328;
        mem[1] = 10'h1d7;
        mem[2] = 10'h1bc;
        mem[3] = 10'h021;
        mem[4] = 10'h240;
        mem[5] = 10'h22e;
        mem[6] = 10'h3c3;
        mem[7] = 10'h188;
        mem[8] = 10'h03a;
        mem[9] = 10'h354;
        mem[10] = 10'h0b4;
        mem[11] = 10'h0f8;
        mem[12] = 10'h1d1;
        mem[13] = 10'h332;
        mem[14] = 10'h09a;
        mem[15] = 10'h132;
        mem[16] = 10'h2a8;
        mem[17] = 10'h080;
        mem[18] = 10'h1ef;
        mem[19] = 10'h12c;
        mem[20] = 10'h166;
        mem[21] = 10'h14a;
        mem[22] = 10'h157;
        mem[23] = 10'h1a5;
        mem[24] = 10'h3d3;
        mem[25] = 10'h24d;
        mem[26] = 10'h23f;
        mem[27] = 10'h3be;
        mem[28] = 10'h2f3;
        mem[29] = 10'h38d;
        mem[30] = 10'h0a3;
        mem[31] = 10'h068;
        mem[32] = 10'h20f;
        mem[33] = 10'h2d5;
        mem[34] = 10'h220;
        mem[35] = 10'h308;
        mem[36] = 10'h3df;
        mem[37] = 10'h0ad;
        mem[38] = 10'h3b1;
        mem[39] = 10'h318;
        mem[40] = 10'h3f6;
        mem[41] = 10'h1f7;
        mem[42] = 10'h0e1;
        mem[43] = 10'h02f;
        mem[44] = 10'h187;
        mem[45] = 10'h29a;
        mem[46] = 10'h195;
        mem[47] = 10'h3c6;
        mem[48] = 10'h2fd;
        mem[49] = 10'h314;
        mem[50] = 10'h03e;
        mem[51] = 10'h172;
        mem[52] = 10'h366;
        mem[53] = 10'h1cf;
        mem[54] = 10'h1ca;
        mem[55] = 10'h317;
        mem[56] = 10'h0e9;
        mem[57] = 10'h324;
        mem[58] = 10'h129;
        mem[59] = 10'h365;
        mem[60] = 10'h38e;
        mem[61] = 10'h1f2;
        mem[62] = 10'h35e;
        mem[63] = 10'h199;
        mem[64] = 10'h2af;
        mem[65] = 10'h3ac;
        mem[66] = 10'h256;
        mem[67] = 10'h06a;
        mem[68] = 10'h34f;
        mem[69] = 10'h1c7;
        mem[70] = 10'h037;
        mem[71] = 10'h21d;
        mem[72] = 10'h311;
        mem[73] = 10'h0ae;
        mem[74] = 10'h15b;
        mem[75] = 10'h3bb;
        mem[76] = 10'h277;
        mem[77] = 10'h338;
        mem[78] = 10'h1c6;
        mem[79] = 10'h33e;
        mem[80] = 10'h25c;
        mem[81] = 10'h171;
        mem[82] = 10'h32f;
        mem[83] = 10'h3da;
        mem[84] = 10'h18f;
        mem[85] = 10'h3d9;
        mem[86] = 10'h08c;
        mem[87] = 10'h0d0;
        mem[88] = 10'h1b2;
        mem[89] = 10'h2e6;
        mem[90] = 10'h159;
        mem[91] = 10'h34b;
        mem[92] = 10'h01b;
        mem[93] = 10'h2c0;
        mem[94] = 10'h020;
        mem[95] = 10'h23c;
        mem[96] = 10'h09f;
        mem[97] = 10'h085;
        mem[98] = 10'h12a;
        mem[99] = 10'h0e7;
        mem[100] = 10'h140;
        mem[101] = 10'h1b0;
        mem[102] = 10'h1b3;
        mem[103] = 10'h185;
        mem[104] = 10'h3a1;
        mem[105] = 10'h051;
        mem[106] = 10'h379;
        mem[107] = 10'h12b;
        mem[108] = 10'h1a0;
        mem[109] = 10'h26e;
        mem[110] = 10'h24e;
        mem[111] = 10'h326;
        mem[112] = 10'h3f0;
        mem[113] = 10'h2ab;
        mem[114] = 10'h35f;
        mem[115] = 10'h1d2;
        mem[116] = 10'h028;
        mem[117] = 10'h3b9;
        mem[118] = 10'h052;
        mem[119] = 10'h078;
        mem[120] = 10'h2f6;
        mem[121] = 10'h3ec;
        mem[122] = 10'h2b2;
        mem[123] = 10'h3f5;
        mem[124] = 10'h226;
        mem[125] = 10'h18b;
        mem[126] = 10'h1bd;
        mem[127] = 10'h0ab;
        mem[128] = 10'h3dd;
        mem[129] = 10'h384;
        mem[130] = 10'h28c;
        mem[131] = 10'h38a;
        mem[132] = 10'h21b;
        mem[133] = 10'h34a;
        mem[134] = 10'h067;
        mem[135] = 10'h180;
        mem[136] = 10'h0a2;
        mem[137] = 10'h170;
        mem[138] = 10'h177;
        mem[139] = 10'h2f1;
        mem[140] = 10'h23b;
        mem[141] = 10'h103;
        mem[142] = 10'h053;
        mem[143] = 10'h3fd;
        mem[144] = 10'h133;
        mem[145] = 10'h275;
        mem[146] = 10'h305;
        mem[147] = 10'h13f;
        mem[148] = 10'h0fa;
        mem[149] = 10'h2d9;
        mem[150] = 10'h29f;
        mem[151] = 10'h2e4;
        mem[152] = 10'h3d7;
        mem[153] = 10'h261;
        mem[154] = 10'h113;
        mem[155] = 10'h230;
        mem[156] = 10'h155;
        mem[157] = 10'h3b5;
        mem[158] = 10'h1f6;
        mem[159] = 10'h22d;
        mem[160] = 10'h386;
        mem[161] = 10'h0dc;
        mem[162] = 10'h0b2;
        mem[163] = 10'h0eb;
        mem[164] = 10'h20a;
        mem[165] = 10'h264;
        mem[166] = 10'h1bf;
        mem[167] = 10'h19e;
        mem[168] = 10'h35a;
        mem[169] = 10'h06e;
        mem[170] = 10'h225;
        mem[171] = 10'h217;
        mem[172] = 10'h3b6;
        mem[173] = 10'h1d5;
        mem[174] = 10'h2b1;
        mem[175] = 10'h055;
        mem[176] = 10'h347;
        mem[177] = 10'h060;
        mem[178] = 10'h3cf;
        mem[179] = 10'h0b7;
        mem[180] = 10'h087;
        mem[181] = 10'h3ff;
        mem[182] = 10'h1f1;
        mem[183] = 10'h156;
        mem[184] = 10'h0d7;
        mem[185] = 10'h197;
        mem[186] = 10'h239;
        mem[187] = 10'h389;
        mem[188] = 10'h1e9;
        mem[189] = 10'h02d;
        mem[190] = 10'h284;
        mem[191] = 10'h145;
        mem[192] = 10'h3d0;
        mem[193] = 10'h375;
        mem[194] = 10'h1ba;
        mem[195] = 10'h331;
        mem[196] = 10'h2ba;
        mem[197] = 10'h07f;
        mem[198] = 10'h20b;
        mem[199] = 10'h254;
        mem[200] = 10'h0d5;
        mem[201] = 10'h0ac;
        mem[202] = 10'h3ca;
        mem[203] = 10'h127;
        mem[204] = 10'h16d;
        mem[205] = 10'h2c6;
        mem[206] = 10'h0a7;
        mem[207] = 10'h0a6;
        mem[208] = 10'h095;
        mem[209] = 10'h179;
        mem[210] = 10'h27d;
        mem[211] = 10'h11c;
        mem[212] = 10'h2f0;
        mem[213] = 10'h16b;
        mem[214] = 10'h0bf;
        mem[215] = 10'h31b;
        mem[216] = 10'h13a;
        mem[217] = 10'h198;
        mem[218] = 10'h320;
        mem[219] = 10'h3bd;
        mem[220] = 10'h0be;
        mem[221] = 10'h25f;
        mem[222] = 10'h161;
        mem[223] = 10'h124;
        mem[224] = 10'h0ed;
        mem[225] = 10'h34c;
        mem[226] = 10'h17d;
        mem[227] = 10'h297;
        mem[228] = 10'h203;
        mem[229] = 10'h3cc;
        mem[230] = 10'h1ee;
        mem[231] = 10'h3c8;
        mem[232] = 10'h2dc;
        mem[233] = 10'h076;
        mem[234] = 10'h094;
        mem[235] = 10'h2ee;
        mem[236] = 10'h265;
        mem[237] = 10'h12d;
        mem[238] = 10'h0b0;
        mem[239] = 10'h205;
        mem[240] = 10'h20d;
        mem[241] = 10'h01d;
        mem[242] = 10'h02c;
        mem[243] = 10'h23e;
        mem[244] = 10'h09e;
        mem[245] = 10'h0d1;
        mem[246] = 10'h353;
        mem[247] = 10'h3bf;
        mem[248] = 10'h089;
        mem[249] = 10'h351;
        mem[250] = 10'h0de;
        mem[251] = 10'h290;
        mem[252] = 10'h06f;
        mem[253] = 10'h00a;
        mem[254] = 10'h0ef;
        mem[255] = 10'h05c;
        mem[256] = 10'h16c;
        mem[257] = 10'h201;
        mem[258] = 10'h36a;
        mem[259] = 10'h1e2;
        mem[260] = 10'h1d6;
        mem[261] = 10'h2d0;
        mem[262] = 10'h015;
        mem[263] = 10'h27a;
        mem[264] = 10'h31e;
        mem[265] = 10'h0ff;
        mem[266] = 10'h3b7;
        mem[267] = 10'h259;
        mem[268] = 10'h3fc;
        mem[269] = 10'h3a7;
        mem[270] = 10'h01c;
        mem[271] = 10'h36f;
        mem[272] = 10'h000;
        mem[273] = 10'h04b;
        mem[274] = 10'h181;
        mem[275] = 10'h0b8;
        mem[276] = 10'h13b;
        mem[277] = 10'h30d;
        mem[278] = 10'h1b1;
        mem[279] = 10'h1a1;
        mem[280] = 10'h05e;
        mem[281] = 10'h21f;
        mem[282] = 10'h126;
        mem[283] = 10'h193;
        mem[284] = 10'h2f5;
        mem[285] = 10'h14c;
        mem[286] = 10'h070;
        mem[287] = 10'h1b6;
        mem[288] = 10'h0c1;
        mem[289] = 10'h35d;
        mem[290] = 10'h0aa;
        mem[291] = 10'h3e1;
        mem[292] = 10'h2d6;
        mem[293] = 10'h19b;
        mem[294] = 10'h13d;
        mem[295] = 10'h144;
        mem[296] = 10'h2e9;
        mem[297] = 10'h1c5;
        mem[298] = 10'h2da;
        mem[299] = 10'h2d7;
        mem[300] = 10'h2cf;
        mem[301] = 10'h003;
        mem[302] = 10'h1f9;
        mem[303] = 10'h056;
        mem[304] = 10'h1cd;
        mem[305] = 10'h1c8;
        mem[306] = 10'h10c;
        mem[307] = 10'h28f;
        mem[308] = 10'h044;
        mem[309] = 10'h380;
        mem[310] = 10'h260;
        mem[311] = 10'h05f;
        mem[312] = 10'h2b7;
        mem[313] = 10'h153;
        mem[314] = 10'h139;
        mem[315] = 10'h345;
        mem[316] = 10'h3b2;
        mem[317] = 10'h1aa;
        mem[318] = 10'h151;
        mem[319] = 10'h300;
        mem[320] = 10'h025;
        mem[321] = 10'h33a;
        mem[322] = 10'h1af;
        mem[323] = 10'h1f3;
        mem[324] = 10'h3a5;
        mem[325] = 10'h3e8;
        mem[326] = 10'h269;
        mem[327] = 10'h105;
        mem[328] = 10'h097;
        mem[329] = 10'h35b;
        mem[330] = 10'h152;
        mem[331] = 10'h0a0;
        mem[332] = 10'h38c;
        mem[333] = 10'h128;
        mem[334] = 10'h271;
        mem[335] = 10'h253;
        mem[336] = 10'h358;
        mem[337] = 10'h3af;
        mem[338] = 10'h2e2;
        mem[339] = 10'h1c9;
        mem[340] = 10'h04f;
        mem[341] = 10'h03b;
        mem[342] = 10'h11d;
        mem[343] = 10'h221;
        mem[344] = 10'h31c;
        mem[345] = 10'h232;
        mem[346] = 10'h32e;
        mem[347] = 10'h1f5;
        mem[348] = 10'h002;
        mem[349] = 10'h377;
        mem[350] = 10'h169;
        mem[351] = 10'h1ad;
        mem[352] = 10'h017;
        mem[353] = 10'h0d4;
        mem[354] = 10'h093;
        mem[355] = 10'h143;
        mem[356] = 10'h285;
        mem[357] = 10'h022;
        mem[358] = 10'h149;
        mem[359] = 10'h17e;
        mem[360] = 10'h21c;
        mem[361] = 10'h2d3;
        mem[362] = 10'h244;
        mem[363] = 10'h245;
        mem[364] = 10'h1cb;
        mem[365] = 10'h3a0;
        mem[366] = 10'h10d;
        mem[367] = 10'h14e;
        mem[368] = 10'h1e5;
        mem[369] = 10'h369;
        mem[370] = 10'h234;
        mem[371] = 10'h372;
        mem[372] = 10'h196;
        mem[373] = 10'h3ed;
        mem[374] = 10'h248;
        mem[375] = 10'h09c;
        mem[376] = 10'h32b;
        mem[377] = 10'h3f2;
        mem[378] = 10'h0f4;
        mem[379] = 10'h2d1;
        mem[380] = 10'h28e;
        mem[381] = 10'h2a7;
        mem[382] = 10'h37e;
        mem[383] = 10'h148;
        mem[384] = 10'h299;
        mem[385] = 10'h267;
        mem[386] = 10'h39a;
        mem[387] = 10'h1e7;
        mem[388] = 10'h0e3;
        mem[389] = 10'h2de;
        mem[390] = 10'h2ac;
        mem[391] = 10'h3c0;
        mem[392] = 10'h363;
        mem[393] = 10'h123;
        mem[394] = 10'h2dd;
        mem[395] = 10'h26b;
        mem[396] = 10'h2ae;
        mem[397] = 10'h235;
        mem[398] = 10'h121;
        mem[399] = 10'h361;
        mem[400] = 10'h323;
        mem[401] = 10'h255;
        mem[402] = 10'h23a;
        mem[403] = 10'h229;
        mem[404] = 10'h0fe;
        mem[405] = 10'h1db;
        mem[406] = 10'h202;
        mem[407] = 10'h288;
        mem[408] = 10'h088;
        mem[409] = 10'h17f;
        mem[410] = 10'h03c;
        mem[411] = 10'h2bd;
        mem[412] = 10'h266;
        mem[413] = 10'h2fe;
        mem[414] = 10'h3bc;
        mem[415] = 10'h2cd;
        mem[416] = 10'h09b;
        mem[417] = 10'h208;
        mem[418] = 10'h31f;
        mem[419] = 10'h399;
        mem[420] = 10'h2d8;
        mem[421] = 10'h15a;
        mem[422] = 10'h340;
        mem[423] = 10'h29b;
        mem[424] = 10'h382;
        mem[425] = 10'h357;
        mem[426] = 10'h390;
        mem[427] = 10'h392;
        mem[428] = 10'h11e;
        mem[429] = 10'h1b4;
        mem[430] = 10'h355;
        mem[431] = 10'h303;
        mem[432] = 10'h039;
        mem[433] = 10'h16a;
        mem[434] = 10'h3fe;
        mem[435] = 10'h310;
        mem[436] = 10'h079;
        mem[437] = 10'h25e;
        mem[438] = 10'h135;
        mem[439] = 10'h316;
        mem[440] = 10'h081;
        mem[441] = 10'h122;
        mem[442] = 10'h33b;
        mem[443] = 10'h295;
        mem[444] = 10'h327;
        mem[445] = 10'h0c0;
        mem[446] = 10'h019;
        mem[447] = 10'h348;
        mem[448] = 10'h05d;
        mem[449] = 10'h05b;
        mem[450] = 10'h2f2;
        mem[451] = 10'h01a;
        mem[452] = 10'h3a3;
        mem[453] = 10'h36e;
        mem[454] = 10'h385;
        mem[455] = 10'h2d2;
        mem[456] = 10'h0c8;
        mem[457] = 10'h370;
        mem[458] = 10'h2e3;
        mem[459] = 10'h1d0;
        mem[460] = 10'h3ef;
        mem[461] = 10'h37b;
        mem[462] = 10'h2cb;
        mem[463] = 10'h24b;
        mem[464] = 10'h114;
        mem[465] = 10'h330;
        mem[466] = 10'h3c5;
        mem[467] = 10'h3a4;
        mem[468] = 10'h0e6;
        mem[469] = 10'h298;
        mem[470] = 10'h045;
        mem[471] = 10'h219;
        mem[472] = 10'h34e;
        mem[473] = 10'h31d;
        mem[474] = 10'h1a7;
        mem[475] = 10'h336;
        mem[476] = 10'h1c1;
        mem[477] = 10'h339;
        mem[478] = 10'h18a;
        mem[479] = 10'h25b;
        mem[480] = 10'h0f7;
        mem[481] = 10'h19d;
        mem[482] = 10'h37a;
        mem[483] = 10'h0b6;
        mem[484] = 10'h191;
        mem[485] = 10'h31a;
        mem[486] = 10'h024;
        mem[487] = 10'h168;
        mem[488] = 10'h342;
        mem[489] = 10'h102;
        mem[490] = 10'h007;
        mem[491] = 10'h138;
        mem[492] = 10'h012;
        mem[493] = 10'h29c;
        mem[494] = 10'h0f3;
        mem[495] = 10'h117;
        mem[496] = 10'h26d;
        mem[497] = 10'h0c5;
        mem[498] = 10'h3f1;
        mem[499] = 10'h341;
        mem[500] = 10'h150;
        mem[501] = 10'h2b0;
        mem[502] = 10'h3c2;
        mem[503] = 10'h32d;
        mem[504] = 10'h061;
        mem[505] = 10'h21e;
        mem[506] = 10'h1fb;
        mem[507] = 10'h218;
        mem[508] = 10'h2ea;
        mem[509] = 10'h2a4;
        mem[510] = 10'h39e;
        mem[511] = 10'h071;
        mem[512] = 10'h02e;
        mem[513] = 10'h005;
        mem[514] = 10'h1f8;
        mem[515] = 10'h3e6;
        mem[516] = 10'h325;
        mem[517] = 10'h0b1;
        mem[518] = 10'h20e;
        mem[519] = 10'h0f1;
        mem[520] = 10'h343;
        mem[521] = 10'h397;
        mem[522] = 10'h083;
        mem[523] = 10'h396;
        mem[524] = 10'h190;
        mem[525] = 10'h356;
        mem[526] = 10'h064;
        mem[527] = 10'h39d;
        mem[528] = 10'h0a9;
        mem[529] = 10'h0e2;
        mem[530] = 10'h2e7;
        mem[531] = 10'h1fd;
        mem[532] = 10'h2f8;
        mem[533] = 10'h066;
        mem[534] = 10'h06c;
        mem[535] = 10'h173;
        mem[536] = 10'h041;
        mem[537] = 10'h23d;
        mem[538] = 10'h359;
        mem[539] = 10'h1da;
        mem[540] = 10'h28a;
        mem[541] = 10'h291;
        mem[542] = 10'h047;
        mem[543] = 10'h049;
        mem[544] = 10'h2bb;
        mem[545] = 10'h04c;
        mem[546] = 10'h24f;
        mem[547] = 10'h19c;
        mem[548] = 10'h2d4;
        mem[549] = 10'h24c;
        mem[550] = 10'h029;
        mem[551] = 10'h2c3;
        mem[552] = 10'h043;
        mem[553] = 10'h337;
        mem[554] = 10'h031;
        mem[555] = 10'h30a;
        mem[556] = 10'h131;
        mem[557] = 10'h1ab;
        mem[558] = 10'h22b;
        mem[559] = 10'h091;
        mem[560] = 10'h2e8;
        mem[561] = 10'h090;
        mem[562] = 10'h0bd;
        mem[563] = 10'h3b8;
        mem[564] = 10'h37f;
        mem[565] = 10'h0cd;
        mem[566] = 10'h222;
        mem[567] = 10'h2cc;
        mem[568] = 10'h213;
        mem[569] = 10'h3a8;
        mem[570] = 10'h0f9;
        mem[571] = 10'h33c;
        mem[572] = 10'h3e9;
        mem[573] = 10'h13e;
        mem[574] = 10'h246;
        mem[575] = 10'h352;
        mem[576] = 10'h184;
        mem[577] = 10'h3d6;
        mem[578] = 10'h3b3;
        mem[579] = 10'h368;
        mem[580] = 10'h00b;
        mem[581] = 10'h272;
        mem[582] = 10'h373;
        mem[583] = 10'h287;
        mem[584] = 10'h27b;
        mem[585] = 10'h034;
        mem[586] = 10'h04e;
        mem[587] = 10'h1bb;
        mem[588] = 10'h206;
        mem[589] = 10'h350;
        mem[590] = 10'h2eb;
        mem[591] = 10'h099;
        mem[592] = 10'h119;
        mem[593] = 10'h334;
        mem[594] = 10'h2c9;
        mem[595] = 10'h1dd;
        mem[596] = 10'h142;
        mem[597] = 10'h073;
        mem[598] = 10'h3c9;
        mem[599] = 10'h2b8;
        mem[600] = 10'h118;
        mem[601] = 10'h0a5;
        mem[602] = 10'h03d;
        mem[603] = 10'h3ae;
        mem[604] = 10'h160;
        mem[605] = 10'h27e;
        mem[606] = 10'h1a4;
        mem[607] = 10'h186;
        mem[608] = 10'h1df;
        mem[609] = 10'h387;
        mem[610] = 10'h011;
        mem[611] = 10'h063;
        mem[612] = 10'h112;
        mem[613] = 10'h10a;
        mem[614] = 10'h06d;
        mem[615] = 10'h293;
        mem[616] = 10'h14d;
        mem[617] = 10'h378;
        mem[618] = 10'h249;
        mem[619] = 10'h141;
        mem[620] = 10'h086;
        mem[621] = 10'h212;
        mem[622] = 10'h302;
        mem[623] = 10'h2be;
        mem[624] = 10'h367;
        mem[625] = 10'h364;
        mem[626] = 10'h042;
        mem[627] = 10'h29e;
        mem[628] = 10'h035;
        mem[629] = 10'h178;
        mem[630] = 10'h1a6;
        mem[631] = 10'h0ba;
        mem[632] = 10'h2c1;
        mem[633] = 10'h39b;
        mem[634] = 10'h074;
        mem[635] = 10'h1d4;
        mem[636] = 10'h1b7;
        mem[637] = 10'h3c7;
        mem[638] = 10'h3fa;
        mem[639] = 10'h2bc;
        mem[640] = 10'h033;
        mem[641] = 10'h0fc;
        mem[642] = 10'h3e4;
        mem[643] = 10'h120;
        mem[644] = 10'h26c;
        mem[645] = 10'h07d;
        mem[646] = 10'h391;
        mem[647] = 10'h15c;
        mem[648] = 10'h2a9;
        mem[649] = 10'h237;
        mem[650] = 10'h3dc;
        mem[651] = 10'h26f;
        mem[652] = 10'h309;
        mem[653] = 10'h100;
        mem[654] = 10'h21a;
        mem[655] = 10'h1a2;
        mem[656] = 10'h16e;
        mem[657] = 10'h010;
        mem[658] = 10'h2b4;
        mem[659] = 10'h3c4;
        mem[660] = 10'h2c2;
        mem[661] = 10'h3f7;
        mem[662] = 10'h1ea;
        mem[663] = 10'h0c2;
        mem[664] = 10'h1e1;
        mem[665] = 10'h3e5;
        mem[666] = 10'h00c;
        mem[667] = 10'h0f6;
        mem[668] = 10'h02b;
        mem[669] = 10'h0c3;
        mem[670] = 10'h2c5;
        mem[671] = 10'h294;
        mem[672] = 10'h3ce;
        mem[673] = 10'h238;
        mem[674] = 10'h3e7;
        mem[675] = 10'h17a;
        mem[676] = 10'h349;
        mem[677] = 10'h242;
        mem[678] = 10'h1eb;
        mem[679] = 10'h136;
        mem[680] = 10'h08e;
        mem[681] = 10'h1fc;
        mem[682] = 10'h2b6;
        mem[683] = 10'h315;
        mem[684] = 10'h00d;
        mem[685] = 10'h147;
        mem[686] = 10'h0bc;
        mem[687] = 10'h28b;
        mem[688] = 10'h39c;
        mem[689] = 10'h09d;
        mem[690] = 10'h1d3;
        mem[691] = 10'h3a6;
        mem[692] = 10'h236;
        mem[693] = 10'h3d5;
        mem[694] = 10'h1fa;
        mem[695] = 10'h281;
        mem[696] = 10'h274;
        mem[697] = 10'h125;
        mem[698] = 10'h3a2;
        mem[699] = 10'h395;
        mem[700] = 10'h069;
        mem[701] = 10'h381;
        mem[702] = 10'h01e;
        mem[703] = 10'h0e0;
        mem[704] = 10'h2a1;
        mem[705] = 10'h233;
        mem[706] = 10'h32a;
        mem[707] = 10'h30e;
        mem[708] = 10'h2a5;
        mem[709] = 10'h2c4;
        mem[710] = 10'h1dc;
        mem[711] = 10'h02a;
        mem[712] = 10'h0cb;
        mem[713] = 10'h106;
        mem[714] = 10'h030;
        mem[715] = 10'h3b0;
        mem[716] = 10'h258;
        mem[717] = 10'h062;
        mem[718] = 10'h279;
        mem[719] = 10'h2e0;
        mem[720] = 10'h174;
        mem[721] = 10'h1d9;
        mem[722] = 10'h250;
        mem[723] = 10'h12e;
        mem[724] = 10'h296;
        mem[725] = 10'h32c;
        mem[726] = 10'h335;
        mem[727] = 10'h1e0;
        mem[728] = 10'h07b;
        mem[729] = 10'h301;
        mem[730] = 10'h360;
        mem[731] = 10'h194;
        mem[732] = 10'h292;
        mem[733] = 10'h398;
        mem[734] = 10'h032;
        mem[735] = 10'h0c9;
        mem[736] = 10'h22c;
        mem[737] = 10'h0cf;
        mem[738] = 10'h0a8;
        mem[739] = 10'h3f8;
        mem[740] = 10'h03f;
        mem[741] = 10'h0d2;
        mem[742] = 10'h215;
        mem[743] = 10'h1e4;
        mem[744] = 10'h2ef;
        mem[745] = 10'h1c0;
        mem[746] = 10'h11a;
        mem[747] = 10'h2f4;
        mem[748] = 10'h065;
        mem[749] = 10'h307;
        mem[750] = 10'h00f;
        mem[751] = 10'h0da;
        mem[752] = 10'h0a4;
        mem[753] = 10'h231;
        mem[754] = 10'h3e0;
        mem[755] = 10'h228;
        mem[756] = 10'h17b;
        mem[757] = 10'h223;
        mem[758] = 10'h06b;
        mem[759] = 10'h3f9;
        mem[760] = 10'h2a2;
        mem[761] = 10'h20c;
        mem[762] = 10'h1e6;
        mem[763] = 10'h1a9;
        mem[764] = 10'h0ca;
        mem[765] = 10'h22a;
        mem[766] = 10'h050;
        mem[767] = 10'h059;
        mem[768] = 10'h077;
        mem[769] = 10'h158;
        mem[770] = 10'h3f4;
        mem[771] = 10'h2ec;
        mem[772] = 10'h25d;
        mem[773] = 10'h0cc;
        mem[774] = 10'h30f;
        mem[775] = 10'h3a9;
        mem[776] = 10'h36c;
        mem[777] = 10'h0df;
        mem[778] = 10'h004;
        mem[779] = 10'h137;
        mem[780] = 10'h006;
        mem[781] = 10'h19a;
        mem[782] = 10'h3aa;
        mem[783] = 10'h29d;
        mem[784] = 10'h276;
        mem[785] = 10'h1a8;
        mem[786] = 10'h04a;
        mem[787] = 10'h3d8;
        mem[788] = 10'h0c4;
        mem[789] = 10'h312;
        mem[790] = 10'h0ce;
        mem[791] = 10'h0fd;
        mem[792] = 10'h1b9;
        mem[793] = 10'h210;
        mem[794] = 10'h18c;
        mem[795] = 10'h3b4;
        mem[796] = 10'h3d2;
        mem[797] = 10'h27c;
        mem[798] = 10'h3eb;
        mem[799] = 10'h263;
        mem[800] = 10'h18d;
        mem[801] = 10'h014;
        mem[802] = 10'h082;
        mem[803] = 10'h075;
        mem[804] = 10'h164;
        mem[805] = 10'h2ad;
        mem[806] = 10'h2ed;
        mem[807] = 10'h36d;
        mem[808] = 10'h108;
        mem[809] = 10'h046;
        mem[810] = 10'h24a;
        mem[811] = 10'h319;
        mem[812] = 10'h34d;
        mem[813] = 10'h0e4;
        mem[814] = 10'h0c6;
        mem[815] = 10'h322;
        mem[816] = 10'h058;
        mem[817] = 10'h0d9;
        mem[818] = 10'h0af;
        mem[819] = 10'h115;
        mem[820] = 10'h1ae;
        mem[821] = 10'h2fa;
        mem[822] = 10'h209;
        mem[823] = 10'h3d1;
        mem[824] = 10'h247;
        mem[825] = 10'h2ca;
        mem[826] = 10'h15e;
        mem[827] = 10'h224;
        mem[828] = 10'h163;
        mem[829] = 10'h252;
        mem[830] = 10'h3cd;
        mem[831] = 10'h1b8;
        mem[832] = 10'h009;
        mem[833] = 10'h008;
        mem[834] = 10'h176;
        mem[835] = 10'h07c;
        mem[836] = 10'h072;
        mem[837] = 10'h040;
        mem[838] = 10'h0c7;
        mem[839] = 10'h2b9;
        mem[840] = 10'h28d;
        mem[841] = 10'h01f;
        mem[842] = 10'h19f;
        mem[843] = 10'h0f0;
        mem[844] = 10'h2c8;
        mem[845] = 10'h251;
        mem[846] = 10'h154;
        mem[847] = 10'h38f;
        mem[848] = 10'h3de;
        mem[849] = 10'h33d;
        mem[850] = 10'h37d;
        mem[851] = 10'h1ec;
        mem[852] = 10'h0f5;
        mem[853] = 10'h27f;
        mem[854] = 10'h2e1;
        mem[855] = 10'h241;
        mem[856] = 10'h2a0;
        mem[857] = 10'h22f;
        mem[858] = 10'h167;
        mem[859] = 10'h023;
        mem[860] = 10'h2f7;
        mem[861] = 10'h204;
        mem[862] = 10'h027;
        mem[863] = 10'h2ff;
        mem[864] = 10'h393;
        mem[865] = 10'h092;
        mem[866] = 10'h2fb;
        mem[867] = 10'h10f;
        mem[868] = 10'h329;
        mem[869] = 10'h313;
        mem[870] = 10'h2a3;
        mem[871] = 10'h346;
        mem[872] = 10'h1be;
        mem[873] = 10'h048;
        mem[874] = 10'h14f;
        mem[875] = 10'h268;
        mem[876] = 10'h1c2;
        mem[877] = 10'h0bb;
        mem[878] = 10'h3c1;
        mem[879] = 10'h1fe;
        mem[880] = 10'h211;
        mem[881] = 10'h096;
        mem[882] = 10'h038;
        mem[883] = 10'h013;
        mem[884] = 10'h162;
        mem[885] = 10'h110;
        mem[886] = 10'h101;
        mem[887] = 10'h07e;
        mem[888] = 10'h17c;
        mem[889] = 10'h2fc;
        mem[890] = 10'h0a1;
        mem[891] = 10'h2b3;
        mem[892] = 10'h306;
        mem[893] = 10'h134;
        mem[894] = 10'h15d;
        mem[895] = 10'h018;
        mem[896] = 10'h25a;
        mem[897] = 10'h109;
        mem[898] = 10'h026;
        mem[899] = 10'h130;
        mem[900] = 10'h2e5;
        mem[901] = 10'h08b;
        mem[902] = 10'h243;
        mem[903] = 10'h30c;
        mem[904] = 10'h37c;
        mem[905] = 10'h175;
        mem[906] = 10'h289;
        mem[907] = 10'h036;
        mem[908] = 10'h304;
        mem[909] = 10'h111;
        mem[910] = 10'h283;
        mem[911] = 10'h14b;
        mem[912] = 10'h371;
        mem[913] = 10'h1a3;
        mem[914] = 10'h13c;
        mem[915] = 10'h1ce;
        mem[916] = 10'h3ad;
        mem[917] = 10'h0b5;
        mem[918] = 10'h3f3;
        mem[919] = 10'h1ff;
        mem[920] = 10'h3db;
        mem[921] = 10'h3ba;
        mem[922] = 10'h1ed;
        mem[923] = 10'h11b;
        mem[924] = 10'h0ee;
        mem[925] = 10'h2db;
        mem[926] = 10'h3ee;
        mem[927] = 10'h278;
        mem[928] = 10'h388;
        mem[929] = 10'h0d8;
        mem[930] = 10'h321;
        mem[931] = 10'h1e8;
        mem[932] = 10'h35c;
        mem[933] = 10'h11f;
        mem[934] = 10'h39f;
        mem[935] = 10'h227;
        mem[936] = 10'h1f4;
        mem[937] = 10'h280;
        mem[938] = 10'h383;
        mem[939] = 10'h3fb;
        mem[940] = 10'h15f;
        mem[941] = 10'h374;
        mem[942] = 10'h26a;
        mem[943] = 10'h0ea;
        mem[944] = 10'h2aa;
        mem[945] = 10'h12f;
        mem[946] = 10'h2b5;
        mem[947] = 10'h394;
        mem[948] = 10'h2c7;
        mem[949] = 10'h107;
        mem[950] = 10'h10b;
        mem[951] = 10'h0f2;
        mem[952] = 10'h273;
        mem[953] = 10'h192;
        mem[954] = 10'h3ab;
        mem[955] = 10'h0ec;
        mem[956] = 10'h0dd;
        mem[957] = 10'h10e;
        mem[958] = 10'h3d4;
        mem[959] = 10'h07a;
        mem[960] = 10'h333;
        mem[961] = 10'h001;
        mem[962] = 10'h146;
        mem[963] = 10'h2ce;
        mem[964] = 10'h016;
        mem[965] = 10'h0b3;
        mem[966] = 10'h0d3;
        mem[967] = 10'h104;
        mem[968] = 10'h084;
        mem[969] = 10'h08f;
        mem[970] = 10'h05a;
        mem[971] = 10'h189;
        mem[972] = 10'h262;
        mem[973] = 10'h38b;
        mem[974] = 10'h057;
        mem[975] = 10'h1ac;
        mem[976] = 10'h2df;
        mem[977] = 10'h362;
        mem[978] = 10'h08a;
        mem[979] = 10'h0fb;
        mem[980] = 10'h2f9;
        mem[981] = 10'h1e3;
        mem[982] = 10'h08d;
        mem[983] = 10'h2a6;
        mem[984] = 10'h282;
        mem[985] = 10'h0db;
        mem[986] = 10'h098;
        mem[987] = 10'h3e2;
        mem[988] = 10'h200;
        mem[989] = 10'h1d8;
        mem[990] = 10'h1c3;
        mem[991] = 10'h116;
        mem[992] = 10'h182;
        mem[993] = 10'h270;
        mem[994] = 10'h1b5;
        mem[995] = 10'h216;
        mem[996] = 10'h344;
        mem[997] = 10'h04d;
        mem[998] = 10'h376;
        mem[999] = 10'h0b9;
        mem[1000] = 10'h214;
        mem[1001] = 10'h0e8;
        mem[1002] = 10'h3cb;
        mem[1003] = 10'h3ea;
        mem[1004] = 10'h33f;
        mem[1005] = 10'h36b;
        mem[1006] = 10'h1c4;
        mem[1007] = 10'h183;
        mem[1008] = 10'h054;
        mem[1009] = 10'h0d6;
        mem[1010] = 10'h0e5;
        mem[1011] = 10'h3e3;
        mem[1012] = 10'h00e;
        mem[1013] = 10'h30b;
        mem[1014] = 10'h257;
        mem[1015] = 10'h2bf;
        mem[1016] = 10'h207;
        mem[1017] = 10'h1cc;
        mem[1018] = 10'h165;
        mem[1019] = 10'h16f;
        mem[1020] = 10'h18e;
        mem[1021] = 10'h1f0;
        mem[1022] = 10'h1de;
        mem[1023] = 10'h286;
    end
endmodule

module odo_sbox_large4(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h0bb;
        mem[1] = 10'h284;
        mem[2] = 10'h1f2;
        mem[3] = 10'h3d4;
        mem[4] = 10'h173;
        mem[5] = 10'h15d;
        mem[6] = 10'h2f2;
        mem[7] = 10'h120;
        mem[8] = 10'h104;
        mem[9] = 10'h057;
        mem[10] = 10'h19a;
        mem[11] = 10'h270;
        mem[12] = 10'h08f;
        mem[13] = 10'h351;
        mem[14] = 10'h009;
        mem[15] = 10'h0f0;
        mem[16] = 10'h096;
        mem[17] = 10'h035;
        mem[18] = 10'h0d0;
        mem[19] = 10'h1da;
        mem[20] = 10'h046;
        mem[21] = 10'h3de;
        mem[22] = 10'h08d;
        mem[23] = 10'h144;
        mem[24] = 10'h148;
        mem[25] = 10'h1a3;
        mem[26] = 10'h164;
        mem[27] = 10'h09f;
        mem[28] = 10'h1d6;
        mem[29] = 10'h3a2;
        mem[30] = 10'h056;
        mem[31] = 10'h0ab;
        mem[32] = 10'h3a6;
        mem[33] = 10'h22e;
        mem[34] = 10'h128;
        mem[35] = 10'h08b;
        mem[36] = 10'h20e;
        mem[37] = 10'h2fa;
        mem[38] = 10'h039;
        mem[39] = 10'h12a;
        mem[40] = 10'h01e;
        mem[41] = 10'h35e;
        mem[42] = 10'h2b4;
        mem[43] = 10'h2eb;
        mem[44] = 10'h2d1;
        mem[45] = 10'h310;
        mem[46] = 10'h281;
        mem[47] = 10'h2d7;
        mem[48] = 10'h30a;
        mem[49] = 10'h35a;
        mem[50] = 10'h306;
        mem[51] = 10'h1b0;
        mem[52] = 10'h354;
        mem[53] = 10'h286;
        mem[54] = 10'h398;
        mem[55] = 10'h2b0;
        mem[56] = 10'h1fc;
        mem[57] = 10'h29c;
        mem[58] = 10'h2d3;
        mem[59] = 10'h27a;
        mem[60] = 10'h05f;
        mem[61] = 10'h04f;
        mem[62] = 10'h2f4;
        mem[63] = 10'h183;
        mem[64] = 10'h041;
        mem[65] = 10'h0be;
        mem[66] = 10'h045;
        mem[67] = 10'h2d8;
        mem[68] = 10'h00b;
        mem[69] = 10'h2a9;
        mem[70] = 10'h001;
        mem[71] = 10'h1a0;
        mem[72] = 10'h0c2;
        mem[73] = 10'h3cb;
        mem[74] = 10'h3b1;
        mem[75] = 10'h269;
        mem[76] = 10'h0c1;
        mem[77] = 10'h3bf;
        mem[78] = 10'h087;
        mem[79] = 10'h1c8;
        mem[80] = 10'h17d;
        mem[81] = 10'h078;
        mem[82] = 10'h1bb;
        mem[83] = 10'h197;
        mem[84] = 10'h027;
        mem[85] = 10'h036;
        mem[86] = 10'h3ac;
        mem[87] = 10'h213;
        mem[88] = 10'h322;
        mem[89] = 10'h3a8;
        mem[90] = 10'h3c1;
        mem[91] = 10'h141;
        mem[92] = 10'h23e;
        mem[93] = 10'h1b5;
        mem[94] = 10'h253;
        mem[95] = 10'h2cb;
        mem[96] = 10'h1e0;
        mem[97] = 10'h3bc;
        mem[98] = 10'h381;
        mem[99] = 10'h2b9;
        mem[100] = 10'h2a3;
        mem[101] = 10'h218;
        mem[102] = 10'h0e9;
        mem[103] = 10'h1f3;
        mem[104] = 10'h06e;
        mem[105] = 10'h010;
        mem[106] = 10'h1ba;
        mem[107] = 10'h063;
        mem[108] = 10'h15c;
        mem[109] = 10'h379;
        mem[110] = 10'h358;
        mem[111] = 10'h25e;
        mem[112] = 10'h1d7;
        mem[113] = 10'h340;
        mem[114] = 10'h3f3;
        mem[115] = 10'h193;
        mem[116] = 10'h1c9;
        mem[117] = 10'h328;
        mem[118] = 10'h292;
        mem[119] = 10'h107;
        mem[120] = 10'h224;
        mem[121] = 10'h198;
        mem[122] = 10'h233;
        mem[123] = 10'h115;
        mem[124] = 10'h326;
        mem[125] = 10'h00d;
        mem[126] = 10'h29a;
        mem[127] = 10'h1db;
        mem[128] = 10'h3c2;
        mem[129] = 10'h305;
        mem[130] = 10'h086;
        mem[131] = 10'h1f8;
        mem[132] = 10'h162;
        mem[133] = 10'h018;
        mem[134] = 10'h36a;
        mem[135] = 10'h0d2;
        mem[136] = 10'h256;
        mem[137] = 10'h30b;
        mem[138] = 10'h0e2;
        mem[139] = 10'h1b9;
        mem[140] = 10'h016;
        mem[141] = 10'h2d0;
        mem[142] = 10'h39b;
        mem[143] = 10'h249;
        mem[144] = 10'h2a5;
        mem[145] = 10'h108;
        mem[146] = 10'h385;
        mem[147] = 10'h1e4;
        mem[148] = 10'h28a;
        mem[149] = 10'h21e;
        mem[150] = 10'h1c5;
        mem[151] = 10'h268;
        mem[152] = 10'h117;
        mem[153] = 10'h012;
        mem[154] = 10'h22c;
        mem[155] = 10'h014;
        mem[156] = 10'h1b8;
        mem[157] = 10'h203;
        mem[158] = 10'h098;
        mem[159] = 10'h026;
        mem[160] = 10'h00f;
        mem[161] = 10'h38b;
        mem[162] = 10'h0b8;
        mem[163] = 10'h105;
        mem[164] = 10'h346;
        mem[165] = 10'h068;
        mem[166] = 10'h075;
        mem[167] = 10'h33e;
        mem[168] = 10'h24c;
        mem[169] = 10'h047;
        mem[170] = 10'h16e;
        mem[171] = 10'h051;
        mem[172] = 10'h0d9;
        mem[173] = 10'h14e;
        mem[174] = 10'h146;
        mem[175] = 10'h2c7;
        mem[176] = 10'h1c7;
        mem[177] = 10'h0ba;
        mem[178] = 10'h24e;
        mem[179] = 10'h2b8;
        mem[180] = 10'h13e;
        mem[181] = 10'h2f5;
        mem[182] = 10'h0c8;
        mem[183] = 10'h19b;
        mem[184] = 10'h327;
        mem[185] = 10'h149;
        mem[186] = 10'h0e5;
        mem[187] = 10'h3d3;
        mem[188] = 10'h366;
        mem[189] = 10'h067;
        mem[190] = 10'h1ce;
        mem[191] = 10'h0f1;
        mem[192] = 10'h2c5;
        mem[193] = 10'h2ae;
        mem[194] = 10'h29e;
        mem[195] = 10'h3b0;
        mem[196] = 10'h3ea;
        mem[197] = 10'h00e;
        mem[198] = 10'h1ec;
        mem[199] = 10'h11b;
        mem[200] = 10'h39e;
        mem[201] = 10'h00a;
        mem[202] = 10'h015;
        mem[203] = 10'h1f9;
        mem[204] = 10'h02e;
        mem[205] = 10'h1df;
        mem[206] = 10'h178;
        mem[207] = 10'h2f1;
        mem[208] = 10'h308;
        mem[209] = 10'h25d;
        mem[210] = 10'h0f3;
        mem[211] = 10'h2f8;
        mem[212] = 10'h1ef;
        mem[213] = 10'h023;
        mem[214] = 10'h1a7;
        mem[215] = 10'h2e5;
        mem[216] = 10'h1e5;
        mem[217] = 10'h1dd;
        mem[218] = 10'h33b;
        mem[219] = 10'h23a;
        mem[220] = 10'h07b;
        mem[221] = 10'h3d0;
        mem[222] = 10'h396;
        mem[223] = 10'h03a;
        mem[224] = 10'h177;
        mem[225] = 10'h3db;
        mem[226] = 10'h368;
        mem[227] = 10'h0e0;
        mem[228] = 10'h35c;
        mem[229] = 10'h196;
        mem[230] = 10'h2b6;
        mem[231] = 10'h1ca;
        mem[232] = 10'h341;
        mem[233] = 10'h0fa;
        mem[234] = 10'h26e;
        mem[235] = 10'h37b;
        mem[236] = 10'h27b;
        mem[237] = 10'h19c;
        mem[238] = 10'h07a;
        mem[239] = 10'h3fe;
        mem[240] = 10'h2cf;
        mem[241] = 10'h37d;
        mem[242] = 10'h034;
        mem[243] = 10'h132;
        mem[244] = 10'h091;
        mem[245] = 10'h3af;
        mem[246] = 10'h0d4;
        mem[247] = 10'h01d;
        mem[248] = 10'h004;
        mem[249] = 10'h158;
        mem[250] = 10'h18f;
        mem[251] = 10'h229;
        mem[252] = 10'h0f2;
        mem[253] = 10'h153;
        mem[254] = 10'h3e7;
        mem[255] = 10'h071;
        mem[256] = 10'h16c;
        mem[257] = 10'h3fc;
        mem[258] = 10'h13f;
        mem[259] = 10'h1e8;
        mem[260] = 10'h3ae;
        mem[261] = 10'h303;
        mem[262] = 10'h2cd;
        mem[263] = 10'h1e2;
        mem[264] = 10'h150;
        mem[265] = 10'h382;
        mem[266] = 10'h3a7;
        mem[267] = 10'h3cf;
        mem[268] = 10'h3e3;
        mem[269] = 10'h013;
        mem[270] = 10'h2aa;
        mem[271] = 10'h099;
        mem[272] = 10'h232;
        mem[273] = 10'h29f;
        mem[274] = 10'h200;
        mem[275] = 10'h113;
        mem[276] = 10'h384;
        mem[277] = 10'h219;
        mem[278] = 10'h126;
        mem[279] = 10'h22d;
        mem[280] = 10'h26c;
        mem[281] = 10'h208;
        mem[282] = 10'h23c;
        mem[283] = 10'h185;
        mem[284] = 10'h1e7;
        mem[285] = 10'h0f7;
        mem[286] = 10'h0c6;
        mem[287] = 10'h102;
        mem[288] = 10'h339;
        mem[289] = 10'h276;
        mem[290] = 10'h09e;
        mem[291] = 10'h2b5;
        mem[292] = 10'h08e;
        mem[293] = 10'h3a5;
        mem[294] = 10'h01b;
        mem[295] = 10'h263;
        mem[296] = 10'h184;
        mem[297] = 10'h1e9;
        mem[298] = 10'h1fd;
        mem[299] = 10'h0ea;
        mem[300] = 10'h1bf;
        mem[301] = 10'h191;
        mem[302] = 10'h138;
        mem[303] = 10'h25b;
        mem[304] = 10'h15b;
        mem[305] = 10'h246;
        mem[306] = 10'h006;
        mem[307] = 10'h2d2;
        mem[308] = 10'h139;
        mem[309] = 10'h2cc;
        mem[310] = 10'h312;
        mem[311] = 10'h3d9;
        mem[312] = 10'h27d;
        mem[313] = 10'h364;
        mem[314] = 10'h255;
        mem[315] = 10'h31e;
        mem[316] = 10'h14d;
        mem[317] = 10'h336;
        mem[318] = 10'h27f;
        mem[319] = 10'h2fc;
        mem[320] = 10'h202;
        mem[321] = 10'h134;
        mem[322] = 10'h282;
        mem[323] = 10'h19e;
        mem[324] = 10'h15a;
        mem[325] = 10'h293;
        mem[326] = 10'h2bc;
        mem[327] = 10'h1e1;
        mem[328] = 10'h337;
        mem[329] = 10'h13a;
        mem[330] = 10'h2d4;
        mem[331] = 10'h1cc;
        mem[332] = 10'h1ee;
        mem[333] = 10'h17a;
        mem[334] = 10'h34e;
        mem[335] = 10'h1e6;
        mem[336] = 10'h3d5;
        mem[337] = 10'h1b6;
        mem[338] = 10'h0b5;
        mem[339] = 10'h359;
        mem[340] = 10'h050;
        mem[341] = 10'h1c4;
        mem[342] = 10'h3cc;
        mem[343] = 10'h301;
        mem[344] = 10'h0f8;
        mem[345] = 10'h302;
        mem[346] = 10'h23f;
        mem[347] = 10'h080;
        mem[348] = 10'h2ff;
        mem[349] = 10'h297;
        mem[350] = 10'h0ff;
        mem[351] = 10'h2a1;
        mem[352] = 10'h168;
        mem[353] = 10'h2b3;
        mem[354] = 10'h028;
        mem[355] = 10'h189;
        mem[356] = 10'h397;
        mem[357] = 10'h0ec;
        mem[358] = 10'h076;
        mem[359] = 10'h058;
        mem[360] = 10'h378;
        mem[361] = 10'h27c;
        mem[362] = 10'h23d;
        mem[363] = 10'h3a4;
        mem[364] = 10'h319;
        mem[365] = 10'h1c0;
        mem[366] = 10'h2a4;
        mem[367] = 10'h3a9;
        mem[368] = 10'h22f;
        mem[369] = 10'h157;
        mem[370] = 10'h3ef;
        mem[371] = 10'h35b;
        mem[372] = 10'h059;
        mem[373] = 10'h331;
        mem[374] = 10'h0cd;
        mem[375] = 10'h257;
        mem[376] = 10'h0cc;
        mem[377] = 10'h12d;
        mem[378] = 10'h2ad;
        mem[379] = 10'h227;
        mem[380] = 10'h2f9;
        mem[381] = 10'h2b2;
        mem[382] = 10'h186;
        mem[383] = 10'h362;
        mem[384] = 10'h2dc;
        mem[385] = 10'h10d;
        mem[386] = 10'h365;
        mem[387] = 10'h3f8;
        mem[388] = 10'h0f9;
        mem[389] = 10'h272;
        mem[390] = 10'h399;
        mem[391] = 10'h205;
        mem[392] = 10'h291;
        mem[393] = 10'h30f;
        mem[394] = 10'h06c;
        mem[395] = 10'h352;
        mem[396] = 10'h350;
        mem[397] = 10'h221;
        mem[398] = 10'h06d;
        mem[399] = 10'h0d8;
        mem[400] = 10'h0eb;
        mem[401] = 10'h357;
        mem[402] = 10'h179;
        mem[403] = 10'h0b0;
        mem[404] = 10'h290;
        mem[405] = 10'h22a;
        mem[406] = 10'h04c;
        mem[407] = 10'h2c1;
        mem[408] = 10'h36c;
        mem[409] = 10'h372;
        mem[410] = 10'h011;
        mem[411] = 10'h055;
        mem[412] = 10'h373;
        mem[413] = 10'h14b;
        mem[414] = 10'h0aa;
        mem[415] = 10'h159;
        mem[416] = 10'h288;
        mem[417] = 10'h040;
        mem[418] = 10'h17e;
        mem[419] = 10'h389;
        mem[420] = 10'h374;
        mem[421] = 10'h020;
        mem[422] = 10'h304;
        mem[423] = 10'h181;
        mem[424] = 10'h3b9;
        mem[425] = 10'h332;
        mem[426] = 10'h033;
        mem[427] = 10'h343;
        mem[428] = 10'h118;
        mem[429] = 10'h31a;
        mem[430] = 10'h0c7;
        mem[431] = 10'h05a;
        mem[432] = 10'h1e3;
        mem[433] = 10'h11f;
        mem[434] = 10'h049;
        mem[435] = 10'h3fb;
        mem[436] = 10'h24d;
        mem[437] = 10'h1af;
        mem[438] = 10'h38c;
        mem[439] = 10'h33c;
        mem[440] = 10'h3ce;
        mem[441] = 10'h147;
        mem[442] = 10'h14a;
        mem[443] = 10'h239;
        mem[444] = 10'h172;
        mem[445] = 10'h05d;
        mem[446] = 10'h3f2;
        mem[447] = 10'h31f;
        mem[448] = 10'h1d3;
        mem[449] = 10'h2f6;
        mem[450] = 10'h21b;
        mem[451] = 10'h3a3;
        mem[452] = 10'h3c7;
        mem[453] = 10'h02c;
        mem[454] = 10'h1fb;
        mem[455] = 10'h02d;
        mem[456] = 10'h022;
        mem[457] = 10'h252;
        mem[458] = 10'h13d;
        mem[459] = 10'h161;
        mem[460] = 10'h28e;
        mem[461] = 10'h2e0;
        mem[462] = 10'h3c9;
        mem[463] = 10'h1dc;
        mem[464] = 10'h390;
        mem[465] = 10'h10e;
        mem[466] = 10'h130;
        mem[467] = 10'h3bd;
        mem[468] = 10'h2c2;
        mem[469] = 10'h1b1;
        mem[470] = 10'h31b;
        mem[471] = 10'h1a2;
        mem[472] = 10'h235;
        mem[473] = 10'h2de;
        mem[474] = 10'h3da;
        mem[475] = 10'h199;
        mem[476] = 10'h26f;
        mem[477] = 10'h38a;
        mem[478] = 10'h29d;
        mem[479] = 10'h3f4;
        mem[480] = 10'h066;
        mem[481] = 10'h002;
        mem[482] = 10'h04b;
        mem[483] = 10'h3d6;
        mem[484] = 10'h36b;
        mem[485] = 10'h261;
        mem[486] = 10'h0fc;
        mem[487] = 10'h182;
        mem[488] = 10'h156;
        mem[489] = 10'h2ef;
        mem[490] = 10'h094;
        mem[491] = 10'h296;
        mem[492] = 10'h12e;
        mem[493] = 10'h0ae;
        mem[494] = 10'h3c5;
        mem[495] = 10'h0b9;
        mem[496] = 10'h000;
        mem[497] = 10'h26d;
        mem[498] = 10'h206;
        mem[499] = 10'h042;
        mem[500] = 10'h3c8;
        mem[501] = 10'h007;
        mem[502] = 10'h114;
        mem[503] = 10'h07e;
        mem[504] = 10'h1ed;
        mem[505] = 10'h29b;
        mem[506] = 10'h39a;
        mem[507] = 10'h103;
        mem[508] = 10'h3d8;
        mem[509] = 10'h021;
        mem[510] = 10'h31d;
        mem[511] = 10'h079;
        mem[512] = 10'h264;
        mem[513] = 10'h0c5;
        mem[514] = 10'h13b;
        mem[515] = 10'h3ad;
        mem[516] = 10'h267;
        mem[517] = 10'h285;
        mem[518] = 10'h122;
        mem[519] = 10'h01f;
        mem[520] = 10'h03f;
        mem[521] = 10'h212;
        mem[522] = 10'h192;
        mem[523] = 10'h3f9;
        mem[524] = 10'h348;
        mem[525] = 10'h17c;
        mem[526] = 10'h1b7;
        mem[527] = 10'h165;
        mem[528] = 10'h34d;
        mem[529] = 10'h25a;
        mem[530] = 10'h031;
        mem[531] = 10'h309;
        mem[532] = 10'h21d;
        mem[533] = 10'h383;
        mem[534] = 10'h258;
        mem[535] = 10'h005;
        mem[536] = 10'h10a;
        mem[537] = 10'h101;
        mem[538] = 10'h060;
        mem[539] = 10'h1cd;
        mem[540] = 10'h2bb;
        mem[541] = 10'h100;
        mem[542] = 10'h215;
        mem[543] = 10'h2a7;
        mem[544] = 10'h3b4;
        mem[545] = 10'h32b;
        mem[546] = 10'h238;
        mem[547] = 10'h1ac;
        mem[548] = 10'h3f7;
        mem[549] = 10'h025;
        mem[550] = 10'h216;
        mem[551] = 10'h345;
        mem[552] = 10'h00c;
        mem[553] = 10'h2a2;
        mem[554] = 10'h24a;
        mem[555] = 10'h2fd;
        mem[556] = 10'h33d;
        mem[557] = 10'h111;
        mem[558] = 10'h0d5;
        mem[559] = 10'h201;
        mem[560] = 10'h2d5;
        mem[561] = 10'h0a7;
        mem[562] = 10'h0dc;
        mem[563] = 10'h0b7;
        mem[564] = 10'h259;
        mem[565] = 10'h0a6;
        mem[566] = 10'h1ae;
        mem[567] = 10'h074;
        mem[568] = 10'h3c3;
        mem[569] = 10'h145;
        mem[570] = 10'h334;
        mem[571] = 10'h20a;
        mem[572] = 10'h3b3;
        mem[573] = 10'h295;
        mem[574] = 10'h1bc;
        mem[575] = 10'h16a;
        mem[576] = 10'h243;
        mem[577] = 10'h0a0;
        mem[578] = 10'h2bf;
        mem[579] = 10'h298;
        mem[580] = 10'h02f;
        mem[581] = 10'h0c0;
        mem[582] = 10'h2be;
        mem[583] = 10'h09d;
        mem[584] = 10'h260;
        mem[585] = 10'h0ee;
        mem[586] = 10'h0fe;
        mem[587] = 10'h323;
        mem[588] = 10'h0e3;
        mem[589] = 10'h3b8;
        mem[590] = 10'h38f;
        mem[591] = 10'h125;
        mem[592] = 10'h376;
        mem[593] = 10'h236;
        mem[594] = 10'h329;
        mem[595] = 10'h1f5;
        mem[596] = 10'h1c2;
        mem[597] = 10'h2a6;
        mem[598] = 10'h017;
        mem[599] = 10'h3ab;
        mem[600] = 10'h38e;
        mem[601] = 10'h28c;
        mem[602] = 10'h1f1;
        mem[603] = 10'h003;
        mem[604] = 10'h1c3;
        mem[605] = 10'h2d6;
        mem[606] = 10'h06a;
        mem[607] = 10'h321;
        mem[608] = 10'h3c6;
        mem[609] = 10'h2ea;
        mem[610] = 10'h084;
        mem[611] = 10'h048;
        mem[612] = 10'h0f4;
        mem[613] = 10'h0bd;
        mem[614] = 10'h053;
        mem[615] = 10'h3f1;
        mem[616] = 10'h28f;
        mem[617] = 10'h195;
        mem[618] = 10'h2e1;
        mem[619] = 10'h18e;
        mem[620] = 10'h2e9;
        mem[621] = 10'h121;
        mem[622] = 10'h36d;
        mem[623] = 10'h277;
        mem[624] = 10'h2b1;
        mem[625] = 10'h01a;
        mem[626] = 10'h054;
        mem[627] = 10'h065;
        mem[628] = 10'h33f;
        mem[629] = 10'h2c8;
        mem[630] = 10'h231;
        mem[631] = 10'h151;
        mem[632] = 10'h265;
        mem[633] = 10'h2db;
        mem[634] = 10'h2df;
        mem[635] = 10'h1de;
        mem[636] = 10'h344;
        mem[637] = 10'h1c6;
        mem[638] = 10'h070;
        mem[639] = 10'h18d;
        mem[640] = 10'h024;
        mem[641] = 10'h38d;
        mem[642] = 10'h3ba;
        mem[643] = 10'h3be;
        mem[644] = 10'h0de;
        mem[645] = 10'h3ff;
        mem[646] = 10'h0fb;
        mem[647] = 10'h24b;
        mem[648] = 10'h10c;
        mem[649] = 10'h388;
        mem[650] = 10'h061;
        mem[651] = 10'h093;
        mem[652] = 10'h247;
        mem[653] = 10'h112;
        mem[654] = 10'h241;
        mem[655] = 10'h211;
        mem[656] = 10'h2ab;
        mem[657] = 10'h1fa;
        mem[658] = 10'h07d;
        mem[659] = 10'h300;
        mem[660] = 10'h3fa;
        mem[661] = 10'h142;
        mem[662] = 10'h20f;
        mem[663] = 10'h380;
        mem[664] = 10'h0e1;
        mem[665] = 10'h0ca;
        mem[666] = 10'h2da;
        mem[667] = 10'h06b;
        mem[668] = 10'h160;
        mem[669] = 10'h3e0;
        mem[670] = 10'h347;
        mem[671] = 10'h089;
        mem[672] = 10'h1ab;
        mem[673] = 10'h273;
        mem[674] = 10'h2ee;
        mem[675] = 10'h03d;
        mem[676] = 10'h2ed;
        mem[677] = 10'h082;
        mem[678] = 10'h25f;
        mem[679] = 10'h1f4;
        mem[680] = 10'h171;
        mem[681] = 10'h029;
        mem[682] = 10'h226;
        mem[683] = 10'h1a9;
        mem[684] = 10'h2c3;
        mem[685] = 10'h0e8;
        mem[686] = 10'h3f0;
        mem[687] = 10'h043;
        mem[688] = 10'h394;
        mem[689] = 10'h3c0;
        mem[690] = 10'h3ee;
        mem[691] = 10'h1d8;
        mem[692] = 10'h03b;
        mem[693] = 10'h170;
        mem[694] = 10'h30c;
        mem[695] = 10'h316;
        mem[696] = 10'h37c;
        mem[697] = 10'h36f;
        mem[698] = 10'h3d7;
        mem[699] = 10'h2c0;
        mem[700] = 10'h0a8;
        mem[701] = 10'h09c;
        mem[702] = 10'h097;
        mem[703] = 10'h0e7;
        mem[704] = 10'h271;
        mem[705] = 10'h393;
        mem[706] = 10'h3e9;
        mem[707] = 10'h129;
        mem[708] = 10'h349;
        mem[709] = 10'h175;
        mem[710] = 10'h0ef;
        mem[711] = 10'h330;
        mem[712] = 10'h180;
        mem[713] = 10'h2fb;
        mem[714] = 10'h2a0;
        mem[715] = 10'h0d1;
        mem[716] = 10'h3d2;
        mem[717] = 10'h05c;
        mem[718] = 10'h15e;
        mem[719] = 10'h05e;
        mem[720] = 10'h392;
        mem[721] = 10'h0b3;
        mem[722] = 10'h395;
        mem[723] = 10'h3c4;
        mem[724] = 10'h3e4;
        mem[725] = 10'h01c;
        mem[726] = 10'h22b;
        mem[727] = 10'h237;
        mem[728] = 10'h3a1;
        mem[729] = 10'h220;
        mem[730] = 10'h275;
        mem[731] = 10'h11d;
        mem[732] = 10'h119;
        mem[733] = 10'h2b7;
        mem[734] = 10'h2ec;
        mem[735] = 10'h2e2;
        mem[736] = 10'h13c;
        mem[737] = 10'h353;
        mem[738] = 10'h3cd;
        mem[739] = 10'h342;
        mem[740] = 10'h0db;
        mem[741] = 10'h131;
        mem[742] = 10'h245;
        mem[743] = 10'h140;
        mem[744] = 10'h315;
        mem[745] = 10'h32f;
        mem[746] = 10'h2e4;
        mem[747] = 10'h0cb;
        mem[748] = 10'h2e8;
        mem[749] = 10'h152;
        mem[750] = 10'h274;
        mem[751] = 10'h3e8;
        mem[752] = 10'h37f;
        mem[753] = 10'h083;
        mem[754] = 10'h325;
        mem[755] = 10'h10f;
        mem[756] = 10'h0f6;
        mem[757] = 10'h2c9;
        mem[758] = 10'h0a3;
        mem[759] = 10'h21c;
        mem[760] = 10'h0a5;
        mem[761] = 10'h11c;
        mem[762] = 10'h044;
        mem[763] = 10'h2dd;
        mem[764] = 10'h2af;
        mem[765] = 10'h39f;
        mem[766] = 10'h210;
        mem[767] = 10'h3ca;
        mem[768] = 10'h0a1;
        mem[769] = 10'h0ce;
        mem[770] = 10'h0c9;
        mem[771] = 10'h167;
        mem[772] = 10'h07c;
        mem[773] = 10'h1eb;
        mem[774] = 10'h135;
        mem[775] = 10'h1a6;
        mem[776] = 10'h222;
        mem[777] = 10'h24f;
        mem[778] = 10'h09a;
        mem[779] = 10'h062;
        mem[780] = 10'h317;
        mem[781] = 10'h02a;
        mem[782] = 10'h3dc;
        mem[783] = 10'h2f3;
        mem[784] = 10'h363;
        mem[785] = 10'h23b;
        mem[786] = 10'h248;
        mem[787] = 10'h223;
        mem[788] = 10'h3f5;
        mem[789] = 10'h1b4;
        mem[790] = 10'h369;
        mem[791] = 10'h1b3;
        mem[792] = 10'h16d;
        mem[793] = 10'h2d9;
        mem[794] = 10'h0c4;
        mem[795] = 10'h110;
        mem[796] = 10'h163;
        mem[797] = 10'h0b2;
        mem[798] = 10'h279;
        mem[799] = 10'h32a;
        mem[800] = 10'h0c3;
        mem[801] = 10'h166;
        mem[802] = 10'h33a;
        mem[803] = 10'h12b;
        mem[804] = 10'h04e;
        mem[805] = 10'h052;
        mem[806] = 10'h31c;
        mem[807] = 10'h0fd;
        mem[808] = 10'h36e;
        mem[809] = 10'h3f6;
        mem[810] = 10'h278;
        mem[811] = 10'h287;
        mem[812] = 10'h1d1;
        mem[813] = 10'h21f;
        mem[814] = 10'h136;
        mem[815] = 10'h0a4;
        mem[816] = 10'h088;
        mem[817] = 10'h04a;
        mem[818] = 10'h11a;
        mem[819] = 10'h1d9;
        mem[820] = 10'h02b;
        mem[821] = 10'h34a;
        mem[822] = 10'h174;
        mem[823] = 10'h037;
        mem[824] = 10'h3d1;
        mem[825] = 10'h1f6;
        mem[826] = 10'h27e;
        mem[827] = 10'h338;
        mem[828] = 10'h09b;
        mem[829] = 10'h371;
        mem[830] = 10'h1be;
        mem[831] = 10'h064;
        mem[832] = 10'h1cf;
        mem[833] = 10'h0ac;
        mem[834] = 10'h214;
        mem[835] = 10'h1ea;
        mem[836] = 10'h3a0;
        mem[837] = 10'h1b2;
        mem[838] = 10'h188;
        mem[839] = 10'h3aa;
        mem[840] = 10'h16f;
        mem[841] = 10'h20d;
        mem[842] = 10'h254;
        mem[843] = 10'h313;
        mem[844] = 10'h1d4;
        mem[845] = 10'h1f7;
        mem[846] = 10'h2c6;
        mem[847] = 10'h1a4;
        mem[848] = 10'h116;
        mem[849] = 10'h3e6;
        mem[850] = 10'h14c;
        mem[851] = 10'h18b;
        mem[852] = 10'h3ec;
        mem[853] = 10'h360;
        mem[854] = 10'h34b;
        mem[855] = 10'h377;
        mem[856] = 10'h032;
        mem[857] = 10'h137;
        mem[858] = 10'h361;
        mem[859] = 10'h39d;
        mem[860] = 10'h250;
        mem[861] = 10'h3dd;
        mem[862] = 10'h21a;
        mem[863] = 10'h0df;
        mem[864] = 10'h240;
        mem[865] = 10'h085;
        mem[866] = 10'h12f;
        mem[867] = 10'h2f0;
        mem[868] = 10'h262;
        mem[869] = 10'h0e6;
        mem[870] = 10'h37e;
        mem[871] = 10'h391;
        mem[872] = 10'h28b;
        mem[873] = 10'h204;
        mem[874] = 10'h18c;
        mem[875] = 10'h244;
        mem[876] = 10'h35f;
        mem[877] = 10'h0b1;
        mem[878] = 10'h283;
        mem[879] = 10'h0e4;
        mem[880] = 10'h127;
        mem[881] = 10'h2ca;
        mem[882] = 10'h324;
        mem[883] = 10'h28d;
        mem[884] = 10'h123;
        mem[885] = 10'h3b6;
        mem[886] = 10'h34f;
        mem[887] = 10'h18a;
        mem[888] = 10'h3b5;
        mem[889] = 10'h375;
        mem[890] = 10'h019;
        mem[891] = 10'h1cb;
        mem[892] = 10'h207;
        mem[893] = 10'h124;
        mem[894] = 10'h1fe;
        mem[895] = 10'h228;
        mem[896] = 10'h370;
        mem[897] = 10'h3e5;
        mem[898] = 10'h038;
        mem[899] = 10'h090;
        mem[900] = 10'h299;
        mem[901] = 10'h1a5;
        mem[902] = 10'h318;
        mem[903] = 10'h2c4;
        mem[904] = 10'h0b6;
        mem[905] = 10'h335;
        mem[906] = 10'h242;
        mem[907] = 10'h0a2;
        mem[908] = 10'h356;
        mem[909] = 10'h0bf;
        mem[910] = 10'h1d0;
        mem[911] = 10'h1c1;
        mem[912] = 10'h17f;
        mem[913] = 10'h2ce;
        mem[914] = 10'h386;
        mem[915] = 10'h26a;
        mem[916] = 10'h367;
        mem[917] = 10'h11e;
        mem[918] = 10'h0d6;
        mem[919] = 10'h187;
        mem[920] = 10'h1aa;
        mem[921] = 10'h34c;
        mem[922] = 10'h307;
        mem[923] = 10'h0cf;
        mem[924] = 10'h10b;
        mem[925] = 10'h32c;
        mem[926] = 10'h0d3;
        mem[927] = 10'h1d5;
        mem[928] = 10'h225;
        mem[929] = 10'h387;
        mem[930] = 10'h081;
        mem[931] = 10'h30e;
        mem[932] = 10'h2fe;
        mem[933] = 10'h3bb;
        mem[934] = 10'h3eb;
        mem[935] = 10'h20b;
        mem[936] = 10'h0a9;
        mem[937] = 10'h095;
        mem[938] = 10'h333;
        mem[939] = 10'h0ad;
        mem[940] = 10'h155;
        mem[941] = 10'h3b7;
        mem[942] = 10'h06f;
        mem[943] = 10'h3ed;
        mem[944] = 10'h143;
        mem[945] = 10'h17b;
        mem[946] = 10'h209;
        mem[947] = 10'h2e7;
        mem[948] = 10'h03e;
        mem[949] = 10'h280;
        mem[950] = 10'h0dd;
        mem[951] = 10'h37a;
        mem[952] = 10'h2ac;
        mem[953] = 10'h16b;
        mem[954] = 10'h20c;
        mem[955] = 10'h355;
        mem[956] = 10'h04d;
        mem[957] = 10'h1d2;
        mem[958] = 10'h19f;
        mem[959] = 10'h092;
        mem[960] = 10'h32e;
        mem[961] = 10'h0da;
        mem[962] = 10'h0f5;
        mem[963] = 10'h154;
        mem[964] = 10'h32d;
        mem[965] = 10'h0bc;
        mem[966] = 10'h08c;
        mem[967] = 10'h07f;
        mem[968] = 10'h25c;
        mem[969] = 10'h3e1;
        mem[970] = 10'h194;
        mem[971] = 10'h190;
        mem[972] = 10'h39c;
        mem[973] = 10'h3e2;
        mem[974] = 10'h2f7;
        mem[975] = 10'h1ff;
        mem[976] = 10'h169;
        mem[977] = 10'h234;
        mem[978] = 10'h1bd;
        mem[979] = 10'h314;
        mem[980] = 10'h251;
        mem[981] = 10'h2e3;
        mem[982] = 10'h0ed;
        mem[983] = 10'h14f;
        mem[984] = 10'h217;
        mem[985] = 10'h12c;
        mem[986] = 10'h133;
        mem[987] = 10'h008;
        mem[988] = 10'h1a1;
        mem[989] = 10'h1f0;
        mem[990] = 10'h289;
        mem[991] = 10'h08a;
        mem[992] = 10'h311;
        mem[993] = 10'h176;
        mem[994] = 10'h03c;
        mem[995] = 10'h05b;
        mem[996] = 10'h077;
        mem[997] = 10'h106;
        mem[998] = 10'h1ad;
        mem[999] = 10'h30d;
        mem[1000] = 10'h35d;
        mem[1001] = 10'h2ba;
        mem[1002] = 10'h072;
        mem[1003] = 10'h3fd;
        mem[1004] = 10'h2a8;
        mem[1005] = 10'h266;
        mem[1006] = 10'h0d7;
        mem[1007] = 10'h3b2;
        mem[1008] = 10'h15f;
        mem[1009] = 10'h294;
        mem[1010] = 10'h2e6;
        mem[1011] = 10'h073;
        mem[1012] = 10'h3df;
        mem[1013] = 10'h230;
        mem[1014] = 10'h030;
        mem[1015] = 10'h1a8;
        mem[1016] = 10'h19d;
        mem[1017] = 10'h069;
        mem[1018] = 10'h0af;
        mem[1019] = 10'h26b;
        mem[1020] = 10'h0b4;
        mem[1021] = 10'h320;
        mem[1022] = 10'h109;
        mem[1023] = 10'h2bd;
    end
endmodule

module odo_sbox_large5(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h103;
        mem[1] = 10'h384;
        mem[2] = 10'h2e6;
        mem[3] = 10'h08c;
        mem[4] = 10'h39d;
        mem[5] = 10'h343;
        mem[6] = 10'h1c5;
        mem[7] = 10'h084;
        mem[8] = 10'h1f0;
        mem[9] = 10'h0a9;
        mem[10] = 10'h2b7;
        mem[11] = 10'h218;
        mem[12] = 10'h1e6;
        mem[13] = 10'h288;
        mem[14] = 10'h3c6;
        mem[15] = 10'h21e;
        mem[16] = 10'h1be;
        mem[17] = 10'h35a;
        mem[18] = 10'h265;
        mem[19] = 10'h118;
        mem[20] = 10'h057;
        mem[21] = 10'h3cb;
        mem[22] = 10'h23e;
        mem[23] = 10'h05a;
        mem[24] = 10'h2da;
        mem[25] = 10'h0aa;
        mem[26] = 10'h128;
        mem[27] = 10'h0c4;
        mem[28] = 10'h352;
        mem[29] = 10'h2c8;
        mem[30] = 10'h0be;
        mem[31] = 10'h3f5;
        mem[32] = 10'h04c;
        mem[33] = 10'h396;
        mem[34] = 10'h195;
        mem[35] = 10'h145;
        mem[36] = 10'h0a5;
        mem[37] = 10'h3f3;
        mem[38] = 10'h1e1;
        mem[39] = 10'h06e;
        mem[40] = 10'h271;
        mem[41] = 10'h108;
        mem[42] = 10'h1c2;
        mem[43] = 10'h19a;
        mem[44] = 10'h2bf;
        mem[45] = 10'h0c8;
        mem[46] = 10'h1ea;
        mem[47] = 10'h309;
        mem[48] = 10'h170;
        mem[49] = 10'h220;
        mem[50] = 10'h1a0;
        mem[51] = 10'h098;
        mem[52] = 10'h125;
        mem[53] = 10'h2bc;
        mem[54] = 10'h12c;
        mem[55] = 10'h2e9;
        mem[56] = 10'h232;
        mem[57] = 10'h03f;
        mem[58] = 10'h0c9;
        mem[59] = 10'h3e3;
        mem[60] = 10'h045;
        mem[61] = 10'h30f;
        mem[62] = 10'h3c7;
        mem[63] = 10'h15b;
        mem[64] = 10'h031;
        mem[65] = 10'h1c8;
        mem[66] = 10'h187;
        mem[67] = 10'h039;
        mem[68] = 10'h04b;
        mem[69] = 10'h101;
        mem[70] = 10'h012;
        mem[71] = 10'h081;
        mem[72] = 10'h139;
        mem[73] = 10'h10f;
        mem[74] = 10'h391;
        mem[75] = 10'h1b9;
        mem[76] = 10'h0a0;
        mem[77] = 10'h2cc;
        mem[78] = 10'h0e9;
        mem[79] = 10'h0de;
        mem[80] = 10'h2ea;
        mem[81] = 10'h33b;
        mem[82] = 10'h191;
        mem[83] = 10'h2c9;
        mem[84] = 10'h3fe;
        mem[85] = 10'h2b5;
        mem[86] = 10'h36e;
        mem[87] = 10'h3a4;
        mem[88] = 10'h397;
        mem[89] = 10'h2c0;
        mem[90] = 10'h3dc;
        mem[91] = 10'h133;
        mem[92] = 10'h252;
        mem[93] = 10'h048;
        mem[94] = 10'h255;
        mem[95] = 10'h33a;
        mem[96] = 10'h0a6;
        mem[97] = 10'h152;
        mem[98] = 10'h149;
        mem[99] = 10'h138;
        mem[100] = 10'h1d1;
        mem[101] = 10'h242;
        mem[102] = 10'h0ec;
        mem[103] = 10'h0ee;
        mem[104] = 10'h003;
        mem[105] = 10'h1fc;
        mem[106] = 10'h2f5;
        mem[107] = 10'h104;
        mem[108] = 10'h39c;
        mem[109] = 10'h0e0;
        mem[110] = 10'h18a;
        mem[111] = 10'h23c;
        mem[112] = 10'h0a3;
        mem[113] = 10'h240;
        mem[114] = 10'h006;
        mem[115] = 10'h03e;
        mem[116] = 10'h12e;
        mem[117] = 10'h338;
        mem[118] = 10'h2df;
        mem[119] = 10'h047;
        mem[120] = 10'h32d;
        mem[121] = 10'h261;
        mem[122] = 10'h2a4;
        mem[123] = 10'h25c;
        mem[124] = 10'h22a;
        mem[125] = 10'h1d9;
        mem[126] = 10'h079;
        mem[127] = 10'h112;
        mem[128] = 10'h3d8;
        mem[129] = 10'h075;
        mem[130] = 10'h221;
        mem[131] = 10'h276;
        mem[132] = 10'h22f;
        mem[133] = 10'h1fb;
        mem[134] = 10'h26a;
        mem[135] = 10'h2c2;
        mem[136] = 10'h1a2;
        mem[137] = 10'h028;
        mem[138] = 10'h07a;
        mem[139] = 10'h353;
        mem[140] = 10'h03b;
        mem[141] = 10'h291;
        mem[142] = 10'h110;
        mem[143] = 10'h1b8;
        mem[144] = 10'h2ba;
        mem[145] = 10'h2c4;
        mem[146] = 10'h284;
        mem[147] = 10'h011;
        mem[148] = 10'h3a8;
        mem[149] = 10'h2cf;
        mem[150] = 10'h08f;
        mem[151] = 10'h364;
        mem[152] = 10'h2d0;
        mem[153] = 10'h026;
        mem[154] = 10'h19f;
        mem[155] = 10'h30e;
        mem[156] = 10'h2f3;
        mem[157] = 10'h2a9;
        mem[158] = 10'h185;
        mem[159] = 10'h222;
        mem[160] = 10'h368;
        mem[161] = 10'h085;
        mem[162] = 10'h09f;
        mem[163] = 10'h1f7;
        mem[164] = 10'h350;
        mem[165] = 10'h31f;
        mem[166] = 10'h1b3;
        mem[167] = 10'h07c;
        mem[168] = 10'h31e;
        mem[169] = 10'h29b;
        mem[170] = 10'h1a7;
        mem[171] = 10'h372;
        mem[172] = 10'h2a8;
        mem[173] = 10'h2f7;
        mem[174] = 10'h229;
        mem[175] = 10'h063;
        mem[176] = 10'h09a;
        mem[177] = 10'h2f1;
        mem[178] = 10'h15a;
        mem[179] = 10'h0b0;
        mem[180] = 10'h0e7;
        mem[181] = 10'h27d;
        mem[182] = 10'h3a2;
        mem[183] = 10'h038;
        mem[184] = 10'h3b5;
        mem[185] = 10'h29c;
        mem[186] = 10'h001;
        mem[187] = 10'h1df;
        mem[188] = 10'h1de;
        mem[189] = 10'h06f;
        mem[190] = 10'h0b2;
        mem[191] = 10'h319;
        mem[192] = 10'h1b6;
        mem[193] = 10'h1d3;
        mem[194] = 10'h3ed;
        mem[195] = 10'h30b;
        mem[196] = 10'h24d;
        mem[197] = 10'h088;
        mem[198] = 10'h3a1;
        mem[199] = 10'h23f;
        mem[200] = 10'h354;
        mem[201] = 10'h27e;
        mem[202] = 10'h245;
        mem[203] = 10'h0ce;
        mem[204] = 10'h377;
        mem[205] = 10'h07f;
        mem[206] = 10'h386;
        mem[207] = 10'h283;
        mem[208] = 10'h0ad;
        mem[209] = 10'h180;
        mem[210] = 10'h11c;
        mem[211] = 10'h13d;
        mem[212] = 10'h019;
        mem[213] = 10'h349;
        mem[214] = 10'h320;
        mem[215] = 10'h080;
        mem[216] = 10'h096;
        mem[217] = 10'h1f3;
        mem[218] = 10'h3d2;
        mem[219] = 10'h325;
        mem[220] = 10'h059;
        mem[221] = 10'h3f7;
        mem[222] = 10'h06a;
        mem[223] = 10'h3b2;
        mem[224] = 10'h0b8;
        mem[225] = 10'h09d;
        mem[226] = 10'h05e;
        mem[227] = 10'h304;
        mem[228] = 10'h1f8;
        mem[229] = 10'h109;
        mem[230] = 10'h3f8;
        mem[231] = 10'h37e;
        mem[232] = 10'h06d;
        mem[233] = 10'h310;
        mem[234] = 10'h280;
        mem[235] = 10'h1a5;
        mem[236] = 10'h3bb;
        mem[237] = 10'h044;
        mem[238] = 10'h34b;
        mem[239] = 10'h077;
        mem[240] = 10'h200;
        mem[241] = 10'h086;
        mem[242] = 10'h04a;
        mem[243] = 10'h18d;
        mem[244] = 10'h127;
        mem[245] = 10'h173;
        mem[246] = 10'h300;
        mem[247] = 10'h296;
        mem[248] = 10'h0dc;
        mem[249] = 10'h398;
        mem[250] = 10'h14f;
        mem[251] = 10'h182;
        mem[252] = 10'h3d7;
        mem[253] = 10'h26b;
        mem[254] = 10'h270;
        mem[255] = 10'h33d;
        mem[256] = 10'h311;
        mem[257] = 10'h3e9;
        mem[258] = 10'h00b;
        mem[259] = 10'h0fe;
        mem[260] = 10'h0eb;
        mem[261] = 10'h0af;
        mem[262] = 10'h32b;
        mem[263] = 10'h093;
        mem[264] = 10'h3fc;
        mem[265] = 10'h0d3;
        mem[266] = 10'h322;
        mem[267] = 10'h022;
        mem[268] = 10'h11e;
        mem[269] = 10'h3a6;
        mem[270] = 10'h3a7;
        mem[271] = 10'h12d;
        mem[272] = 10'h030;
        mem[273] = 10'h263;
        mem[274] = 10'h1c4;
        mem[275] = 10'h068;
        mem[276] = 10'h2b6;
        mem[277] = 10'h226;
        mem[278] = 10'h27a;
        mem[279] = 10'h20a;
        mem[280] = 10'h335;
        mem[281] = 10'h231;
        mem[282] = 10'h326;
        mem[283] = 10'h22e;
        mem[284] = 10'h3e1;
        mem[285] = 10'h16b;
        mem[286] = 10'h137;
        mem[287] = 10'h04f;
        mem[288] = 10'h215;
        mem[289] = 10'h143;
        mem[290] = 10'h33e;
        mem[291] = 10'h2a3;
        mem[292] = 10'h237;
        mem[293] = 10'h367;
        mem[294] = 10'h018;
        mem[295] = 10'h1a4;
        mem[296] = 10'h31c;
        mem[297] = 10'h07b;
        mem[298] = 10'h142;
        mem[299] = 10'h285;
        mem[300] = 10'h09e;
        mem[301] = 10'h100;
        mem[302] = 10'h22b;
        mem[303] = 10'h2b9;
        mem[304] = 10'h040;
        mem[305] = 10'h3ef;
        mem[306] = 10'h1b7;
        mem[307] = 10'h36a;
        mem[308] = 10'h28c;
        mem[309] = 10'h107;
        mem[310] = 10'h28a;
        mem[311] = 10'h2e8;
        mem[312] = 10'h184;
        mem[313] = 10'h0dd;
        mem[314] = 10'h12a;
        mem[315] = 10'h0bf;
        mem[316] = 10'h3d3;
        mem[317] = 10'h3bf;
        mem[318] = 10'h3a3;
        mem[319] = 10'h32e;
        mem[320] = 10'h399;
        mem[321] = 10'h0f7;
        mem[322] = 10'h105;
        mem[323] = 10'h3b4;
        mem[324] = 10'h14b;
        mem[325] = 10'h122;
        mem[326] = 10'h3c8;
        mem[327] = 10'h0bd;
        mem[328] = 10'h15d;
        mem[329] = 10'h01d;
        mem[330] = 10'h095;
        mem[331] = 10'h334;
        mem[332] = 10'h157;
        mem[333] = 10'h3a5;
        mem[334] = 10'h2c5;
        mem[335] = 10'h17a;
        mem[336] = 10'h0e4;
        mem[337] = 10'h192;
        mem[338] = 10'h156;
        mem[339] = 10'h10a;
        mem[340] = 10'h166;
        mem[341] = 10'h094;
        mem[342] = 10'h321;
        mem[343] = 10'h204;
        mem[344] = 10'h00e;
        mem[345] = 10'h1cd;
        mem[346] = 10'h35d;
        mem[347] = 10'h360;
        mem[348] = 10'h297;
        mem[349] = 10'h2f4;
        mem[350] = 10'h37a;
        mem[351] = 10'h2de;
        mem[352] = 10'h268;
        mem[353] = 10'h1a8;
        mem[354] = 10'h2b4;
        mem[355] = 10'h0ae;
        mem[356] = 10'h017;
        mem[357] = 10'h35f;
        mem[358] = 10'h196;
        mem[359] = 10'h3ad;
        mem[360] = 10'h239;
        mem[361] = 10'h235;
        mem[362] = 10'h1bb;
        mem[363] = 10'h0a8;
        mem[364] = 10'h35b;
        mem[365] = 10'h3d5;
        mem[366] = 10'h25f;
        mem[367] = 10'h206;
        mem[368] = 10'h0a7;
        mem[369] = 10'h264;
        mem[370] = 10'h37d;
        mem[371] = 10'h31a;
        mem[372] = 10'h193;
        mem[373] = 10'h0b4;
        mem[374] = 10'h163;
        mem[375] = 10'h070;
        mem[376] = 10'h17b;
        mem[377] = 10'h277;
        mem[378] = 10'h020;
        mem[379] = 10'h0c5;
        mem[380] = 10'h35c;
        mem[381] = 10'h36c;
        mem[382] = 10'h11b;
        mem[383] = 10'h015;
        mem[384] = 10'h38d;
        mem[385] = 10'h3ff;
        mem[386] = 10'h021;
        mem[387] = 10'h0ab;
        mem[388] = 10'h295;
        mem[389] = 10'h2f0;
        mem[390] = 10'h362;
        mem[391] = 10'h340;
        mem[392] = 10'h043;
        mem[393] = 10'h298;
        mem[394] = 10'h1da;
        mem[395] = 10'h0fc;
        mem[396] = 10'h344;
        mem[397] = 10'h302;
        mem[398] = 10'h3f9;
        mem[399] = 10'h1cf;
        mem[400] = 10'h2ab;
        mem[401] = 10'h15e;
        mem[402] = 10'h257;
        mem[403] = 10'h0b5;
        mem[404] = 10'h17e;
        mem[405] = 10'h253;
        mem[406] = 10'h1c0;
        mem[407] = 10'h22c;
        mem[408] = 10'h0ba;
        mem[409] = 10'h36d;
        mem[410] = 10'h275;
        mem[411] = 10'h0f2;
        mem[412] = 10'h3b1;
        mem[413] = 10'h056;
        mem[414] = 10'h3e0;
        mem[415] = 10'h014;
        mem[416] = 10'h119;
        mem[417] = 10'h178;
        mem[418] = 10'h294;
        mem[419] = 10'h3e7;
        mem[420] = 10'h13f;
        mem[421] = 10'h3cf;
        mem[422] = 10'h379;
        mem[423] = 10'h2e2;
        mem[424] = 10'h3b7;
        mem[425] = 10'h3f1;
        mem[426] = 10'h005;
        mem[427] = 10'h008;
        mem[428] = 10'h18c;
        mem[429] = 10'h066;
        mem[430] = 10'h0fa;
        mem[431] = 10'h1af;
        mem[432] = 10'h3ac;
        mem[433] = 10'h342;
        mem[434] = 10'h2b0;
        mem[435] = 10'h301;
        mem[436] = 10'h380;
        mem[437] = 10'h25b;
        mem[438] = 10'h27f;
        mem[439] = 10'h286;
        mem[440] = 10'h383;
        mem[441] = 10'h258;
        mem[442] = 10'h111;
        mem[443] = 10'h02e;
        mem[444] = 10'h331;
        mem[445] = 10'h28e;
        mem[446] = 10'h2f2;
        mem[447] = 10'h256;
        mem[448] = 10'h31d;
        mem[449] = 10'h2a0;
        mem[450] = 10'h176;
        mem[451] = 10'h089;
        mem[452] = 10'h21f;
        mem[453] = 10'h371;
        mem[454] = 10'h3d0;
        mem[455] = 10'h272;
        mem[456] = 10'h1a9;
        mem[457] = 10'h042;
        mem[458] = 10'h14d;
        mem[459] = 10'h1c3;
        mem[460] = 10'h05b;
        mem[461] = 10'h24b;
        mem[462] = 10'h2b1;
        mem[463] = 10'h2d8;
        mem[464] = 10'h22d;
        mem[465] = 10'h369;
        mem[466] = 10'h330;
        mem[467] = 10'h097;
        mem[468] = 10'h073;
        mem[469] = 10'h161;
        mem[470] = 10'h38e;
        mem[471] = 10'h029;
        mem[472] = 10'h027;
        mem[473] = 10'h0d5;
        mem[474] = 10'h062;
        mem[475] = 10'h211;
        mem[476] = 10'h099;
        mem[477] = 10'h058;
        mem[478] = 10'h305;
        mem[479] = 10'h1a1;
        mem[480] = 10'h1e3;
        mem[481] = 10'h1f9;
        mem[482] = 10'h090;
        mem[483] = 10'h385;
        mem[484] = 10'h179;
        mem[485] = 10'h2bb;
        mem[486] = 10'h024;
        mem[487] = 10'h1ab;
        mem[488] = 10'h13a;
        mem[489] = 10'h154;
        mem[490] = 10'h126;
        mem[491] = 10'h370;
        mem[492] = 10'h303;
        mem[493] = 10'h210;
        mem[494] = 10'h21b;
        mem[495] = 10'h1e8;
        mem[496] = 10'h0cf;
        mem[497] = 10'h373;
        mem[498] = 10'h1aa;
        mem[499] = 10'h273;
        mem[500] = 10'h3cd;
        mem[501] = 10'h18f;
        mem[502] = 10'h214;
        mem[503] = 10'h1b4;
        mem[504] = 10'h08d;
        mem[505] = 10'h013;
        mem[506] = 10'h106;
        mem[507] = 10'h316;
        mem[508] = 10'h3a9;
        mem[509] = 10'h17f;
        mem[510] = 10'h1fa;
        mem[511] = 10'h357;
        mem[512] = 10'h19c;
        mem[513] = 10'h3d4;
        mem[514] = 10'h2dd;
        mem[515] = 10'h0c6;
        mem[516] = 10'h217;
        mem[517] = 10'h395;
        mem[518] = 10'h207;
        mem[519] = 10'h3e2;
        mem[520] = 10'h117;
        mem[521] = 10'h3c4;
        mem[522] = 10'h1d0;
        mem[523] = 10'h250;
        mem[524] = 10'h050;
        mem[525] = 10'h26d;
        mem[526] = 10'h1c1;
        mem[527] = 10'h28b;
        mem[528] = 10'h375;
        mem[529] = 10'h060;
        mem[530] = 10'h046;
        mem[531] = 10'h0e6;
        mem[532] = 10'h3aa;
        mem[533] = 10'h293;
        mem[534] = 10'h216;
        mem[535] = 10'h0f9;
        mem[536] = 10'h032;
        mem[537] = 10'h38f;
        mem[538] = 10'h3d1;
        mem[539] = 10'h11d;
        mem[540] = 10'h1b2;
        mem[541] = 10'h121;
        mem[542] = 10'h0c0;
        mem[543] = 10'h25e;
        mem[544] = 10'h189;
        mem[545] = 10'h31b;
        mem[546] = 10'h1e0;
        mem[547] = 10'h2c3;
        mem[548] = 10'h00a;
        mem[549] = 10'h3dd;
        mem[550] = 10'h2f6;
        mem[551] = 10'h3fa;
        mem[552] = 10'h0d1;
        mem[553] = 10'h0ed;
        mem[554] = 10'h212;
        mem[555] = 10'h2a1;
        mem[556] = 10'h11a;
        mem[557] = 10'h0e1;
        mem[558] = 10'h290;
        mem[559] = 10'h3f4;
        mem[560] = 10'h172;
        mem[561] = 10'h205;
        mem[562] = 10'h054;
        mem[563] = 10'h09b;
        mem[564] = 10'h34d;
        mem[565] = 10'h3ae;
        mem[566] = 10'h1f4;
        mem[567] = 10'h287;
        mem[568] = 10'h1e9;
        mem[569] = 10'h233;
        mem[570] = 10'h3f6;
        mem[571] = 10'h091;
        mem[572] = 10'h279;
        mem[573] = 10'h067;
        mem[574] = 10'h129;
        mem[575] = 10'h055;
        mem[576] = 10'h2b3;
        mem[577] = 10'h2eb;
        mem[578] = 10'h36f;
        mem[579] = 10'h1c6;
        mem[580] = 10'h2cd;
        mem[581] = 10'h2ac;
        mem[582] = 10'h14e;
        mem[583] = 10'h16a;
        mem[584] = 10'h382;
        mem[585] = 10'h0a1;
        mem[586] = 10'h289;
        mem[587] = 10'h246;
        mem[588] = 10'h3fb;
        mem[589] = 10'h02c;
        mem[590] = 10'h1b0;
        mem[591] = 10'h356;
        mem[592] = 10'h148;
        mem[593] = 10'h144;
        mem[594] = 10'h2aa;
        mem[595] = 10'h34c;
        mem[596] = 10'h38c;
        mem[597] = 10'h033;
        mem[598] = 10'h315;
        mem[599] = 10'h07d;
        mem[600] = 10'h3b3;
        mem[601] = 10'h1a3;
        mem[602] = 10'h27b;
        mem[603] = 10'h16e;
        mem[604] = 10'h3fd;
        mem[605] = 10'h0cc;
        mem[606] = 10'h113;
        mem[607] = 10'h135;
        mem[608] = 10'h10c;
        mem[609] = 10'h169;
        mem[610] = 10'h333;
        mem[611] = 10'h1d6;
        mem[612] = 10'h238;
        mem[613] = 10'h124;
        mem[614] = 10'h132;
        mem[615] = 10'h1e2;
        mem[616] = 10'h1cc;
        mem[617] = 10'h1d5;
        mem[618] = 10'h3af;
        mem[619] = 10'h0d9;
        mem[620] = 10'h0f1;
        mem[621] = 10'h08e;
        mem[622] = 10'h378;
        mem[623] = 10'h3ea;
        mem[624] = 10'h3ca;
        mem[625] = 10'h102;
        mem[626] = 10'h3ab;
        mem[627] = 10'h38b;
        mem[628] = 10'h376;
        mem[629] = 10'h188;
        mem[630] = 10'h12b;
        mem[631] = 10'h158;
        mem[632] = 10'h36b;
        mem[633] = 10'h09c;
        mem[634] = 10'h136;
        mem[635] = 10'h147;
        mem[636] = 10'h20b;
        mem[637] = 10'h393;
        mem[638] = 10'h2c7;
        mem[639] = 10'h2ad;
        mem[640] = 10'h208;
        mem[641] = 10'h2dc;
        mem[642] = 10'h199;
        mem[643] = 10'h1d8;
        mem[644] = 10'h072;
        mem[645] = 10'h02f;
        mem[646] = 10'h1f6;
        mem[647] = 10'h230;
        mem[648] = 10'h2a5;
        mem[649] = 10'h225;
        mem[650] = 10'h3f2;
        mem[651] = 10'h21a;
        mem[652] = 10'h37f;
        mem[653] = 10'h2a6;
        mem[654] = 10'h1bf;
        mem[655] = 10'h052;
        mem[656] = 10'h1ba;
        mem[657] = 10'h2c6;
        mem[658] = 10'h30d;
        mem[659] = 10'h332;
        mem[660] = 10'h016;
        mem[661] = 10'h0b7;
        mem[662] = 10'h244;
        mem[663] = 10'h2d9;
        mem[664] = 10'h2af;
        mem[665] = 10'h0d6;
        mem[666] = 10'h2ef;
        mem[667] = 10'h313;
        mem[668] = 10'h02d;
        mem[669] = 10'h3c2;
        mem[670] = 10'h05d;
        mem[671] = 10'h282;
        mem[672] = 10'h2d1;
        mem[673] = 10'h19e;
        mem[674] = 10'h1fd;
        mem[675] = 10'h34a;
        mem[676] = 10'h2ae;
        mem[677] = 10'h0ef;
        mem[678] = 10'h04e;
        mem[679] = 10'h308;
        mem[680] = 10'h18b;
        mem[681] = 10'h115;
        mem[682] = 10'h3c0;
        mem[683] = 10'h19d;
        mem[684] = 10'h351;
        mem[685] = 10'h306;
        mem[686] = 10'h17d;
        mem[687] = 10'h0f5;
        mem[688] = 10'h3e8;
        mem[689] = 10'h0a2;
        mem[690] = 10'h00c;
        mem[691] = 10'h361;
        mem[692] = 10'h141;
        mem[693] = 10'h0da;
        mem[694] = 10'h2be;
        mem[695] = 10'h3bc;
        mem[696] = 10'h312;
        mem[697] = 10'h314;
        mem[698] = 10'h15c;
        mem[699] = 10'h39f;
        mem[700] = 10'h3eb;
        mem[701] = 10'h002;
        mem[702] = 10'h3c5;
        mem[703] = 10'h328;
        mem[704] = 10'h0c1;
        mem[705] = 10'h2e0;
        mem[706] = 10'h186;
        mem[707] = 10'h2d3;
        mem[708] = 10'h1ed;
        mem[709] = 10'h0ea;
        mem[710] = 10'h155;
        mem[711] = 10'h25d;
        mem[712] = 10'h247;
        mem[713] = 10'h1e7;
        mem[714] = 10'h1b5;
        mem[715] = 10'h08a;
        mem[716] = 10'h146;
        mem[717] = 10'h0fb;
        mem[718] = 10'h3ce;
        mem[719] = 10'h3ba;
        mem[720] = 10'h174;
        mem[721] = 10'h168;
        mem[722] = 10'h01e;
        mem[723] = 10'h123;
        mem[724] = 10'h0c2;
        mem[725] = 10'h004;
        mem[726] = 10'h0c3;
        mem[727] = 10'h164;
        mem[728] = 10'h387;
        mem[729] = 10'h381;
        mem[730] = 10'h19b;
        mem[731] = 10'h2d4;
        mem[732] = 10'h1c7;
        mem[733] = 10'h1bc;
        mem[734] = 10'h01f;
        mem[735] = 10'h2e4;
        mem[736] = 10'h02a;
        mem[737] = 10'h069;
        mem[738] = 10'h26e;
        mem[739] = 10'h278;
        mem[740] = 10'h14c;
        mem[741] = 10'h114;
        mem[742] = 10'h1f2;
        mem[743] = 10'h3b0;
        mem[744] = 10'h33f;
        mem[745] = 10'h23a;
        mem[746] = 10'h1d2;
        mem[747] = 10'h3d9;
        mem[748] = 10'h010;
        mem[749] = 10'h1c9;
        mem[750] = 10'h336;
        mem[751] = 10'h37b;
        mem[752] = 10'h05c;
        mem[753] = 10'h078;
        mem[754] = 10'h3ec;
        mem[755] = 10'h134;
        mem[756] = 10'h2d7;
        mem[757] = 10'h236;
        mem[758] = 10'h259;
        mem[759] = 10'h227;
        mem[760] = 10'h037;
        mem[761] = 10'h17c;
        mem[762] = 10'h11f;
        mem[763] = 10'h071;
        mem[764] = 10'h162;
        mem[765] = 10'h234;
        mem[766] = 10'h3e4;
        mem[767] = 10'h1e4;
        mem[768] = 10'h0ff;
        mem[769] = 10'h30a;
        mem[770] = 10'h3de;
        mem[771] = 10'h2ff;
        mem[772] = 10'h18e;
        mem[773] = 10'h34e;
        mem[774] = 10'h065;
        mem[775] = 10'h16c;
        mem[776] = 10'h346;
        mem[777] = 10'h12f;
        mem[778] = 10'h249;
        mem[779] = 10'h00f;
        mem[780] = 10'h266;
        mem[781] = 10'h26f;
        mem[782] = 10'h051;
        mem[783] = 10'h2fd;
        mem[784] = 10'h035;
        mem[785] = 10'h0f3;
        mem[786] = 10'h3e6;
        mem[787] = 10'h28d;
        mem[788] = 10'h32f;
        mem[789] = 10'h327;
        mem[790] = 10'h181;
        mem[791] = 10'h116;
        mem[792] = 10'h165;
        mem[793] = 10'h0b6;
        mem[794] = 10'h0c7;
        mem[795] = 10'h05f;
        mem[796] = 10'h0f6;
        mem[797] = 10'h08b;
        mem[798] = 10'h347;
        mem[799] = 10'h1f1;
        mem[800] = 10'h1ad;
        mem[801] = 10'h26c;
        mem[802] = 10'h190;
        mem[803] = 10'h243;
        mem[804] = 10'h2ca;
        mem[805] = 10'h241;
        mem[806] = 10'h281;
        mem[807] = 10'h087;
        mem[808] = 10'h203;
        mem[809] = 10'h0ca;
        mem[810] = 10'h1d4;
        mem[811] = 10'h29f;
        mem[812] = 10'h167;
        mem[813] = 10'h1b1;
        mem[814] = 10'h197;
        mem[815] = 10'h20f;
        mem[816] = 10'h38a;
        mem[817] = 10'h1a6;
        mem[818] = 10'h318;
        mem[819] = 10'h323;
        mem[820] = 10'h339;
        mem[821] = 10'h3b8;
        mem[822] = 10'h0d2;
        mem[823] = 10'h2fb;
        mem[824] = 10'h1ce;
        mem[825] = 10'h2ed;
        mem[826] = 10'h2d2;
        mem[827] = 10'h061;
        mem[828] = 10'h37c;
        mem[829] = 10'h24f;
        mem[830] = 10'h1db;
        mem[831] = 10'h1dc;
        mem[832] = 10'h120;
        mem[833] = 10'h24e;
        mem[834] = 10'h29d;
        mem[835] = 10'h082;
        mem[836] = 10'h1ff;
        mem[837] = 10'h16f;
        mem[838] = 10'h219;
        mem[839] = 10'h317;
        mem[840] = 10'h262;
        mem[841] = 10'h355;
        mem[842] = 10'h0cd;
        mem[843] = 10'h151;
        mem[844] = 10'h3db;
        mem[845] = 10'h32c;
        mem[846] = 10'h0e8;
        mem[847] = 10'h254;
        mem[848] = 10'h269;
        mem[849] = 10'h198;
        mem[850] = 10'h1ca;
        mem[851] = 10'h076;
        mem[852] = 10'h348;
        mem[853] = 10'h159;
        mem[854] = 10'h223;
        mem[855] = 10'h2fa;
        mem[856] = 10'h025;
        mem[857] = 10'h023;
        mem[858] = 10'h2e5;
        mem[859] = 10'h20c;
        mem[860] = 10'h13e;
        mem[861] = 10'h03d;
        mem[862] = 10'h0e2;
        mem[863] = 10'h251;
        mem[864] = 10'h20e;
        mem[865] = 10'h27c;
        mem[866] = 10'h1ae;
        mem[867] = 10'h175;
        mem[868] = 10'h036;
        mem[869] = 10'h213;
        mem[870] = 10'h1bd;
        mem[871] = 10'h130;
        mem[872] = 10'h392;
        mem[873] = 10'h3da;
        mem[874] = 10'h007;
        mem[875] = 10'h1ef;
        mem[876] = 10'h0bb;
        mem[877] = 10'h14a;
        mem[878] = 10'h053;
        mem[879] = 10'h1cb;
        mem[880] = 10'h0f0;
        mem[881] = 10'h329;
        mem[882] = 10'h0e3;
        mem[883] = 10'h194;
        mem[884] = 10'h3b6;
        mem[885] = 10'h01c;
        mem[886] = 10'h292;
        mem[887] = 10'h01b;
        mem[888] = 10'h2a7;
        mem[889] = 10'h25a;
        mem[890] = 10'h13b;
        mem[891] = 10'h2f8;
        mem[892] = 10'h337;
        mem[893] = 10'h201;
        mem[894] = 10'h2fc;
        mem[895] = 10'h0f4;
        mem[896] = 10'h21d;
        mem[897] = 10'h224;
        mem[898] = 10'h3df;
        mem[899] = 10'h1e5;
        mem[900] = 10'h150;
        mem[901] = 10'h1ec;
        mem[902] = 10'h183;
        mem[903] = 10'h32a;
        mem[904] = 10'h0d7;
        mem[905] = 10'h3b9;
        mem[906] = 10'h2e7;
        mem[907] = 10'h06b;
        mem[908] = 10'h35e;
        mem[909] = 10'h0bc;
        mem[910] = 10'h3cc;
        mem[911] = 10'h374;
        mem[912] = 10'h0d8;
        mem[913] = 10'h2a2;
        mem[914] = 10'h083;
        mem[915] = 10'h3d6;
        mem[916] = 10'h3c9;
        mem[917] = 10'h07e;
        mem[918] = 10'h2ce;
        mem[919] = 10'h23d;
        mem[920] = 10'h0b1;
        mem[921] = 10'h2e1;
        mem[922] = 10'h092;
        mem[923] = 10'h04d;
        mem[924] = 10'h0d0;
        mem[925] = 10'h01a;
        mem[926] = 10'h341;
        mem[927] = 10'h29e;
        mem[928] = 10'h1f5;
        mem[929] = 10'h0b9;
        mem[930] = 10'h140;
        mem[931] = 10'h1eb;
        mem[932] = 10'h24a;
        mem[933] = 10'h13c;
        mem[934] = 10'h28f;
        mem[935] = 10'h10e;
        mem[936] = 10'h0fd;
        mem[937] = 10'h00d;
        mem[938] = 10'h0cb;
        mem[939] = 10'h3bd;
        mem[940] = 10'h131;
        mem[941] = 10'h3c3;
        mem[942] = 10'h034;
        mem[943] = 10'h21c;
        mem[944] = 10'h03c;
        mem[945] = 10'h0b3;
        mem[946] = 10'h049;
        mem[947] = 10'h39b;
        mem[948] = 10'h23b;
        mem[949] = 10'h274;
        mem[950] = 10'h33c;
        mem[951] = 10'h228;
        mem[952] = 10'h2c1;
        mem[953] = 10'h359;
        mem[954] = 10'h3a0;
        mem[955] = 10'h02b;
        mem[956] = 10'h390;
        mem[957] = 10'h24c;
        mem[958] = 10'h2cb;
        mem[959] = 10'h10d;
        mem[960] = 10'h0db;
        mem[961] = 10'h1d7;
        mem[962] = 10'h1ac;
        mem[963] = 10'h39e;
        mem[964] = 10'h2b2;
        mem[965] = 10'h202;
        mem[966] = 10'h2e3;
        mem[967] = 10'h160;
        mem[968] = 10'h2ec;
        mem[969] = 10'h16d;
        mem[970] = 10'h2bd;
        mem[971] = 10'h389;
        mem[972] = 10'h39a;
        mem[973] = 10'h074;
        mem[974] = 10'h34f;
        mem[975] = 10'h177;
        mem[976] = 10'h2fe;
        mem[977] = 10'h20d;
        mem[978] = 10'h30c;
        mem[979] = 10'h2f9;
        mem[980] = 10'h10b;
        mem[981] = 10'h363;
        mem[982] = 10'h307;
        mem[983] = 10'h2db;
        mem[984] = 10'h3ee;
        mem[985] = 10'h000;
        mem[986] = 10'h1dd;
        mem[987] = 10'h064;
        mem[988] = 10'h171;
        mem[989] = 10'h2d5;
        mem[990] = 10'h06c;
        mem[991] = 10'h358;
        mem[992] = 10'h3f0;
        mem[993] = 10'h345;
        mem[994] = 10'h0d4;
        mem[995] = 10'h209;
        mem[996] = 10'h1fe;
        mem[997] = 10'h3e5;
        mem[998] = 10'h1ee;
        mem[999] = 10'h03a;
        mem[1000] = 10'h388;
        mem[1001] = 10'h394;
        mem[1002] = 10'h365;
        mem[1003] = 10'h041;
        mem[1004] = 10'h366;
        mem[1005] = 10'h0ac;
        mem[1006] = 10'h0f8;
        mem[1007] = 10'h009;
        mem[1008] = 10'h15f;
        mem[1009] = 10'h299;
        mem[1010] = 10'h2d6;
        mem[1011] = 10'h324;
        mem[1012] = 10'h260;
        mem[1013] = 10'h2ee;
        mem[1014] = 10'h0df;
        mem[1015] = 10'h0e5;
        mem[1016] = 10'h0a4;
        mem[1017] = 10'h2b8;
        mem[1018] = 10'h3c1;
        mem[1019] = 10'h267;
        mem[1020] = 10'h153;
        mem[1021] = 10'h29a;
        mem[1022] = 10'h3be;
        mem[1023] = 10'h248;
    end
endmodule

module odo_sbox_large6(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h185;
        mem[1] = 10'h15e;
        mem[2] = 10'h1a7;
        mem[3] = 10'h0f1;
        mem[4] = 10'h3a2;
        mem[5] = 10'h0e1;
        mem[6] = 10'h18e;
        mem[7] = 10'h2f4;
        mem[8] = 10'h22d;
        mem[9] = 10'h168;
        mem[10] = 10'h3fb;
        mem[11] = 10'h30c;
        mem[12] = 10'h2db;
        mem[13] = 10'h01a;
        mem[14] = 10'h324;
        mem[15] = 10'h0bf;
        mem[16] = 10'h262;
        mem[17] = 10'h348;
        mem[18] = 10'h176;
        mem[19] = 10'h2a8;
        mem[20] = 10'h2d8;
        mem[21] = 10'h1f2;
        mem[22] = 10'h164;
        mem[23] = 10'h3a5;
        mem[24] = 10'h25f;
        mem[25] = 10'h252;
        mem[26] = 10'h307;
        mem[27] = 10'h1d7;
        mem[28] = 10'h3de;
        mem[29] = 10'h219;
        mem[30] = 10'h205;
        mem[31] = 10'h2ef;
        mem[32] = 10'h267;
        mem[33] = 10'h05c;
        mem[34] = 10'h08b;
        mem[35] = 10'h210;
        mem[36] = 10'h1ee;
        mem[37] = 10'h1a2;
        mem[38] = 10'h298;
        mem[39] = 10'h102;
        mem[40] = 10'h0be;
        mem[41] = 10'h3dc;
        mem[42] = 10'h315;
        mem[43] = 10'h195;
        mem[44] = 10'h132;
        mem[45] = 10'h03b;
        mem[46] = 10'h29f;
        mem[47] = 10'h19a;
        mem[48] = 10'h2d1;
        mem[49] = 10'h3a0;
        mem[50] = 10'h3c1;
        mem[51] = 10'h01e;
        mem[52] = 10'h3e7;
        mem[53] = 10'h194;
        mem[54] = 10'h2df;
        mem[55] = 10'h33a;
        mem[56] = 10'h287;
        mem[57] = 10'h29b;
        mem[58] = 10'h116;
        mem[59] = 10'h2af;
        mem[60] = 10'h0af;
        mem[61] = 10'h345;
        mem[62] = 10'h0d1;
        mem[63] = 10'h0ea;
        mem[64] = 10'h3b7;
        mem[65] = 10'h0b8;
        mem[66] = 10'h16d;
        mem[67] = 10'h24e;
        mem[68] = 10'h37a;
        mem[69] = 10'h386;
        mem[70] = 10'h0ff;
        mem[71] = 10'h1b2;
        mem[72] = 10'h1f7;
        mem[73] = 10'h1c4;
        mem[74] = 10'h024;
        mem[75] = 10'h103;
        mem[76] = 10'h001;
        mem[77] = 10'h3d0;
        mem[78] = 10'h20e;
        mem[79] = 10'h26d;
        mem[80] = 10'h099;
        mem[81] = 10'h3fe;
        mem[82] = 10'h1e3;
        mem[83] = 10'h35d;
        mem[84] = 10'h036;
        mem[85] = 10'h23c;
        mem[86] = 10'h1f6;
        mem[87] = 10'h393;
        mem[88] = 10'h0cc;
        mem[89] = 10'h112;
        mem[90] = 10'h3a1;
        mem[91] = 10'h392;
        mem[92] = 10'h041;
        mem[93] = 10'h18b;
        mem[94] = 10'h216;
        mem[95] = 10'h085;
        mem[96] = 10'h22b;
        mem[97] = 10'h0e0;
        mem[98] = 10'h3f5;
        mem[99] = 10'h329;
        mem[100] = 10'h2ba;
        mem[101] = 10'h357;
        mem[102] = 10'h10f;
        mem[103] = 10'h043;
        mem[104] = 10'h117;
        mem[105] = 10'h3a4;
        mem[106] = 10'h30e;
        mem[107] = 10'h07e;
        mem[108] = 10'h359;
        mem[109] = 10'h3e9;
        mem[110] = 10'h2e4;
        mem[111] = 10'h20c;
        mem[112] = 10'h2ee;
        mem[113] = 10'h302;
        mem[114] = 10'h004;
        mem[115] = 10'h0c3;
        mem[116] = 10'h0a4;
        mem[117] = 10'h3f1;
        mem[118] = 10'h1cf;
        mem[119] = 10'h034;
        mem[120] = 10'h032;
        mem[121] = 10'h229;
        mem[122] = 10'h362;
        mem[123] = 10'h05b;
        mem[124] = 10'h15c;
        mem[125] = 10'h3db;
        mem[126] = 10'h276;
        mem[127] = 10'h19b;
        mem[128] = 10'h2a1;
        mem[129] = 10'h0da;
        mem[130] = 10'h27f;
        mem[131] = 10'h1b5;
        mem[132] = 10'h1eb;
        mem[133] = 10'h342;
        mem[134] = 10'h0f9;
        mem[135] = 10'h240;
        mem[136] = 10'h12c;
        mem[137] = 10'h39e;
        mem[138] = 10'h0d3;
        mem[139] = 10'h34d;
        mem[140] = 10'h18d;
        mem[141] = 10'h2c4;
        mem[142] = 10'h1ab;
        mem[143] = 10'h047;
        mem[144] = 10'h3ef;
        mem[145] = 10'h373;
        mem[146] = 10'h361;
        mem[147] = 10'h11e;
        mem[148] = 10'h285;
        mem[149] = 10'h221;
        mem[150] = 10'h2dc;
        mem[151] = 10'h220;
        mem[152] = 10'h217;
        mem[153] = 10'h2e7;
        mem[154] = 10'h0ec;
        mem[155] = 10'h2c7;
        mem[156] = 10'h3f6;
        mem[157] = 10'h069;
        mem[158] = 10'h009;
        mem[159] = 10'h25b;
        mem[160] = 10'h0e3;
        mem[161] = 10'h2a2;
        mem[162] = 10'h0dd;
        mem[163] = 10'h1d5;
        mem[164] = 10'h3b2;
        mem[165] = 10'h376;
        mem[166] = 10'h10d;
        mem[167] = 10'h128;
        mem[168] = 10'h1f5;
        mem[169] = 10'h145;
        mem[170] = 10'h2e1;
        mem[171] = 10'h305;
        mem[172] = 10'h0b4;
        mem[173] = 10'h34a;
        mem[174] = 10'h1fd;
        mem[175] = 10'h388;
        mem[176] = 10'h02e;
        mem[177] = 10'h3b9;
        mem[178] = 10'h390;
        mem[179] = 10'h23d;
        mem[180] = 10'h002;
        mem[181] = 10'h1d6;
        mem[182] = 10'h2a5;
        mem[183] = 10'h1a8;
        mem[184] = 10'h2bb;
        mem[185] = 10'h31f;
        mem[186] = 10'h111;
        mem[187] = 10'h273;
        mem[188] = 10'h2fa;
        mem[189] = 10'h387;
        mem[190] = 10'h17d;
        mem[191] = 10'h3cd;
        mem[192] = 10'h119;
        mem[193] = 10'h02d;
        mem[194] = 10'h044;
        mem[195] = 10'h343;
        mem[196] = 10'h228;
        mem[197] = 10'h0c2;
        mem[198] = 10'h163;
        mem[199] = 10'h148;
        mem[200] = 10'h297;
        mem[201] = 10'h120;
        mem[202] = 10'h0b0;
        mem[203] = 10'h077;
        mem[204] = 10'h1f0;
        mem[205] = 10'h27b;
        mem[206] = 10'h1c9;
        mem[207] = 10'h12d;
        mem[208] = 10'h314;
        mem[209] = 10'h180;
        mem[210] = 10'h2c5;
        mem[211] = 10'h2e6;
        mem[212] = 10'h26e;
        mem[213] = 10'h071;
        mem[214] = 10'h3bd;
        mem[215] = 10'h2b1;
        mem[216] = 10'h1f9;
        mem[217] = 10'h3c6;
        mem[218] = 10'h332;
        mem[219] = 10'h36e;
        mem[220] = 10'h049;
        mem[221] = 10'h06b;
        mem[222] = 10'h0cd;
        mem[223] = 10'h1e9;
        mem[224] = 10'h00e;
        mem[225] = 10'h160;
        mem[226] = 10'h162;
        mem[227] = 10'h126;
        mem[228] = 10'h37e;
        mem[229] = 10'h395;
        mem[230] = 10'h212;
        mem[231] = 10'h3f8;
        mem[232] = 10'h37b;
        mem[233] = 10'h320;
        mem[234] = 10'h33b;
        mem[235] = 10'h123;
        mem[236] = 10'h0df;
        mem[237] = 10'h340;
        mem[238] = 10'h0fb;
        mem[239] = 10'h2e3;
        mem[240] = 10'h1be;
        mem[241] = 10'h0a7;
        mem[242] = 10'h1e2;
        mem[243] = 10'h035;
        mem[244] = 10'h198;
        mem[245] = 10'h17c;
        mem[246] = 10'h26c;
        mem[247] = 10'h31d;
        mem[248] = 10'h32f;
        mem[249] = 10'h23e;
        mem[250] = 10'h28b;
        mem[251] = 10'h060;
        mem[252] = 10'h105;
        mem[253] = 10'h36f;
        mem[254] = 10'h170;
        mem[255] = 10'h0ae;
        mem[256] = 10'h186;
        mem[257] = 10'h309;
        mem[258] = 10'h19e;
        mem[259] = 10'h3ee;
        mem[260] = 10'h149;
        mem[261] = 10'h0a5;
        mem[262] = 10'h19f;
        mem[263] = 10'h183;
        mem[264] = 10'h066;
        mem[265] = 10'h1da;
        mem[266] = 10'h336;
        mem[267] = 10'h0d0;
        mem[268] = 10'h0d8;
        mem[269] = 10'h37d;
        mem[270] = 10'h134;
        mem[271] = 10'h3c0;
        mem[272] = 10'h3d8;
        mem[273] = 10'h057;
        mem[274] = 10'h29a;
        mem[275] = 10'h04d;
        mem[276] = 10'h268;
        mem[277] = 10'h26a;
        mem[278] = 10'h2ec;
        mem[279] = 10'h207;
        mem[280] = 10'h076;
        mem[281] = 10'h1fa;
        mem[282] = 10'h0fc;
        mem[283] = 10'h2d7;
        mem[284] = 10'h21e;
        mem[285] = 10'h1e4;
        mem[286] = 10'h3cc;
        mem[287] = 10'h1f1;
        mem[288] = 10'h274;
        mem[289] = 10'h2dd;
        mem[290] = 10'h21d;
        mem[291] = 10'h265;
        mem[292] = 10'h169;
        mem[293] = 10'h3c7;
        mem[294] = 10'h0d5;
        mem[295] = 10'h09c;
        mem[296] = 10'h3c2;
        mem[297] = 10'h206;
        mem[298] = 10'h22e;
        mem[299] = 10'h211;
        mem[300] = 10'h299;
        mem[301] = 10'h16c;
        mem[302] = 10'h0c4;
        mem[303] = 10'h1e0;
        mem[304] = 10'h003;
        mem[305] = 10'h3e6;
        mem[306] = 10'h28d;
        mem[307] = 10'h04a;
        mem[308] = 10'h25c;
        mem[309] = 10'h073;
        mem[310] = 10'h2de;
        mem[311] = 10'h0cf;
        mem[312] = 10'h1de;
        mem[313] = 10'h3ea;
        mem[314] = 10'h0d4;
        mem[315] = 10'h09b;
        mem[316] = 10'h01b;
        mem[317] = 10'h147;
        mem[318] = 10'h05a;
        mem[319] = 10'h241;
        mem[320] = 10'h3f3;
        mem[321] = 10'h0fe;
        mem[322] = 10'h3e2;
        mem[323] = 10'h0f2;
        mem[324] = 10'h052;
        mem[325] = 10'h3c3;
        mem[326] = 10'h366;
        mem[327] = 10'h033;
        mem[328] = 10'h3c5;
        mem[329] = 10'h18f;
        mem[330] = 10'h3f9;
        mem[331] = 10'h2b2;
        mem[332] = 10'h22c;
        mem[333] = 10'h29c;
        mem[334] = 10'h397;
        mem[335] = 10'h131;
        mem[336] = 10'h0c0;
        mem[337] = 10'h34f;
        mem[338] = 10'h191;
        mem[339] = 10'h20f;
        mem[340] = 10'h013;
        mem[341] = 10'h14e;
        mem[342] = 10'h155;
        mem[343] = 10'h0eb;
        mem[344] = 10'h380;
        mem[345] = 10'h15d;
        mem[346] = 10'h152;
        mem[347] = 10'h25e;
        mem[348] = 10'h21f;
        mem[349] = 10'h050;
        mem[350] = 10'h063;
        mem[351] = 10'h062;
        mem[352] = 10'h233;
        mem[353] = 10'h1c6;
        mem[354] = 10'h172;
        mem[355] = 10'h039;
        mem[356] = 10'h2da;
        mem[357] = 10'h234;
        mem[358] = 10'h264;
        mem[359] = 10'h2bd;
        mem[360] = 10'h254;
        mem[361] = 10'h3ba;
        mem[362] = 10'h322;
        mem[363] = 10'h1f3;
        mem[364] = 10'h215;
        mem[365] = 10'h235;
        mem[366] = 10'h3ae;
        mem[367] = 10'h16f;
        mem[368] = 10'h225;
        mem[369] = 10'h31b;
        mem[370] = 10'h2f5;
        mem[371] = 10'h1df;
        mem[372] = 10'h296;
        mem[373] = 10'h341;
        mem[374] = 10'h243;
        mem[375] = 10'h218;
        mem[376] = 10'h059;
        mem[377] = 10'h025;
        mem[378] = 10'h1bf;
        mem[379] = 10'h2cf;
        mem[380] = 10'h38f;
        mem[381] = 10'h09e;
        mem[382] = 10'h01c;
        mem[383] = 10'h16e;
        mem[384] = 10'h166;
        mem[385] = 10'h09d;
        mem[386] = 10'h2a3;
        mem[387] = 10'h368;
        mem[388] = 10'h01f;
        mem[389] = 10'h1a1;
        mem[390] = 10'h141;
        mem[391] = 10'h095;
        mem[392] = 10'h39f;
        mem[393] = 10'h352;
        mem[394] = 10'h2fe;
        mem[395] = 10'h350;
        mem[396] = 10'h270;
        mem[397] = 10'h21b;
        mem[398] = 10'h3ff;
        mem[399] = 10'h289;
        mem[400] = 10'h0bd;
        mem[401] = 10'h056;
        mem[402] = 10'h203;
        mem[403] = 10'h34e;
        mem[404] = 10'h1e8;
        mem[405] = 10'h28e;
        mem[406] = 10'h091;
        mem[407] = 10'h288;
        mem[408] = 10'h379;
        mem[409] = 10'h2c0;
        mem[410] = 10'h3e1;
        mem[411] = 10'h26f;
        mem[412] = 10'h0c8;
        mem[413] = 10'h150;
        mem[414] = 10'h12f;
        mem[415] = 10'h2f7;
        mem[416] = 10'h1aa;
        mem[417] = 10'h2f6;
        mem[418] = 10'h2b0;
        mem[419] = 10'h2aa;
        mem[420] = 10'h2b4;
        mem[421] = 10'h1ba;
        mem[422] = 10'h3a3;
        mem[423] = 10'h35c;
        mem[424] = 10'h04f;
        mem[425] = 10'h14f;
        mem[426] = 10'h3a9;
        mem[427] = 10'h0e2;
        mem[428] = 10'h0c9;
        mem[429] = 10'h255;
        mem[430] = 10'h08d;
        mem[431] = 10'h23f;
        mem[432] = 10'h37c;
        mem[433] = 10'h0d2;
        mem[434] = 10'h263;
        mem[435] = 10'h171;
        mem[436] = 10'h17e;
        mem[437] = 10'h1b0;
        mem[438] = 10'h2ae;
        mem[439] = 10'h1cc;
        mem[440] = 10'h344;
        mem[441] = 10'h143;
        mem[442] = 10'h281;
        mem[443] = 10'h14c;
        mem[444] = 10'h3e0;
        mem[445] = 10'h382;
        mem[446] = 10'h07a;
        mem[447] = 10'h3d9;
        mem[448] = 10'h101;
        mem[449] = 10'h03d;
        mem[450] = 10'h192;
        mem[451] = 10'h081;
        mem[452] = 10'h3af;
        mem[453] = 10'h2d2;
        mem[454] = 10'h364;
        mem[455] = 10'h1b9;
        mem[456] = 10'h0fa;
        mem[457] = 10'h313;
        mem[458] = 10'h3ac;
        mem[459] = 10'h3ce;
        mem[460] = 10'h29d;
        mem[461] = 10'h040;
        mem[462] = 10'h14b;
        mem[463] = 10'h337;
        mem[464] = 10'h054;
        mem[465] = 10'h136;
        mem[466] = 10'h214;
        mem[467] = 10'h1a3;
        mem[468] = 10'h15b;
        mem[469] = 10'h0b5;
        mem[470] = 10'h027;
        mem[471] = 10'h29e;
        mem[472] = 10'h38a;
        mem[473] = 10'h03e;
        mem[474] = 10'h31a;
        mem[475] = 10'h208;
        mem[476] = 10'h137;
        mem[477] = 10'h3d7;
        mem[478] = 10'h39a;
        mem[479] = 10'h092;
        mem[480] = 10'h000;
        mem[481] = 10'h1c5;
        mem[482] = 10'h083;
        mem[483] = 10'h2eb;
        mem[484] = 10'h399;
        mem[485] = 10'h016;
        mem[486] = 10'h260;
        mem[487] = 10'h0e6;
        mem[488] = 10'h007;
        mem[489] = 10'h38b;
        mem[490] = 10'h283;
        mem[491] = 10'h1ca;
        mem[492] = 10'h292;
        mem[493] = 10'h248;
        mem[494] = 10'h0f5;
        mem[495] = 10'h15a;
        mem[496] = 10'h005;
        mem[497] = 10'h2a6;
        mem[498] = 10'h0a9;
        mem[499] = 10'h202;
        mem[500] = 10'h12a;
        mem[501] = 10'h230;
        mem[502] = 10'h10c;
        mem[503] = 10'h18c;
        mem[504] = 10'h06f;
        mem[505] = 10'h23b;
        mem[506] = 10'h2c8;
        mem[507] = 10'h13a;
        mem[508] = 10'h0a6;
        mem[509] = 10'h279;
        mem[510] = 10'h03c;
        mem[511] = 10'h266;
        mem[512] = 10'h2c2;
        mem[513] = 10'h32b;
        mem[514] = 10'h114;
        mem[515] = 10'h291;
        mem[516] = 10'h097;
        mem[517] = 10'h1ad;
        mem[518] = 10'h086;
        mem[519] = 10'h3e5;
        mem[520] = 10'h03f;
        mem[521] = 10'h1ae;
        mem[522] = 10'h10e;
        mem[523] = 10'h022;
        mem[524] = 10'h261;
        mem[525] = 10'h2ca;
        mem[526] = 10'h25a;
        mem[527] = 10'h072;
        mem[528] = 10'h250;
        mem[529] = 10'h36a;
        mem[530] = 10'h0f3;
        mem[531] = 10'h308;
        mem[532] = 10'h00a;
        mem[533] = 10'h015;
        mem[534] = 10'h3f7;
        mem[535] = 10'h161;
        mem[536] = 10'h2d9;
        mem[537] = 10'h068;
        mem[538] = 10'h1c7;
        mem[539] = 10'h108;
        mem[540] = 10'h061;
        mem[541] = 10'h35a;
        mem[542] = 10'h11c;
        mem[543] = 10'h0ba;
        mem[544] = 10'h2a0;
        mem[545] = 10'h06e;
        mem[546] = 10'h330;
        mem[547] = 10'h3a7;
        mem[548] = 10'h0e5;
        mem[549] = 10'h146;
        mem[550] = 10'h383;
        mem[551] = 10'h316;
        mem[552] = 10'h258;
        mem[553] = 10'h144;
        mem[554] = 10'h100;
        mem[555] = 10'h037;
        mem[556] = 10'h0e4;
        mem[557] = 10'h0b1;
        mem[558] = 10'h360;
        mem[559] = 10'h065;
        mem[560] = 10'h177;
        mem[561] = 10'h242;
        mem[562] = 10'h190;
        mem[563] = 10'h031;
        mem[564] = 10'h30a;
        mem[565] = 10'h1d3;
        mem[566] = 10'h089;
        mem[567] = 10'h27c;
        mem[568] = 10'h3ca;
        mem[569] = 10'h339;
        mem[570] = 10'h12b;
        mem[571] = 10'h2d6;
        mem[572] = 10'h0f0;
        mem[573] = 10'h3dd;
        mem[574] = 10'h1c8;
        mem[575] = 10'h354;
        mem[576] = 10'h07c;
        mem[577] = 10'h338;
        mem[578] = 10'h3d6;
        mem[579] = 10'h37f;
        mem[580] = 10'h21a;
        mem[581] = 10'h385;
        mem[582] = 10'h0ca;
        mem[583] = 10'h30d;
        mem[584] = 10'h2cc;
        mem[585] = 10'h269;
        mem[586] = 10'h334;
        mem[587] = 10'h0ac;
        mem[588] = 10'h1ea;
        mem[589] = 10'h184;
        mem[590] = 10'h3b3;
        mem[591] = 10'h2cb;
        mem[592] = 10'h39c;
        mem[593] = 10'h249;
        mem[594] = 10'h11b;
        mem[595] = 10'h0c6;
        mem[596] = 10'h006;
        mem[597] = 10'h331;
        mem[598] = 10'h2bc;
        mem[599] = 10'h2e9;
        mem[600] = 10'h084;
        mem[601] = 10'h0b6;
        mem[602] = 10'h277;
        mem[603] = 10'h1cb;
        mem[604] = 10'h2c3;
        mem[605] = 10'h13c;
        mem[606] = 10'h33c;
        mem[607] = 10'h226;
        mem[608] = 10'h3fd;
        mem[609] = 10'h067;
        mem[610] = 10'h115;
        mem[611] = 10'h293;
        mem[612] = 10'h1d9;
        mem[613] = 10'h246;
        mem[614] = 10'h0ab;
        mem[615] = 10'h282;
        mem[616] = 10'h32a;
        mem[617] = 10'h1e1;
        mem[618] = 10'h154;
        mem[619] = 10'h303;
        mem[620] = 10'h2d5;
        mem[621] = 10'h353;
        mem[622] = 10'h1b7;
        mem[623] = 10'h17a;
        mem[624] = 10'h2d0;
        mem[625] = 10'h0a3;
        mem[626] = 10'h323;
        mem[627] = 10'h156;
        mem[628] = 10'h369;
        mem[629] = 10'h16a;
        mem[630] = 10'h10b;
        mem[631] = 10'h0e9;
        mem[632] = 10'h023;
        mem[633] = 10'h284;
        mem[634] = 10'h0b3;
        mem[635] = 10'h200;
        mem[636] = 10'h15f;
        mem[637] = 10'h1e6;
        mem[638] = 10'h0ef;
        mem[639] = 10'h370;
        mem[640] = 10'h04b;
        mem[641] = 10'h110;
        mem[642] = 10'h2b8;
        mem[643] = 10'h0d7;
        mem[644] = 10'h028;
        mem[645] = 10'h3fa;
        mem[646] = 10'h1d1;
        mem[647] = 10'h19c;
        mem[648] = 10'h06d;
        mem[649] = 10'h0b7;
        mem[650] = 10'h30b;
        mem[651] = 10'h197;
        mem[652] = 10'h00f;
        mem[653] = 10'h3aa;
        mem[654] = 10'h20b;
        mem[655] = 10'h239;
        mem[656] = 10'h2a7;
        mem[657] = 10'h0f6;
        mem[658] = 10'h107;
        mem[659] = 10'h227;
        mem[660] = 10'h0dc;
        mem[661] = 10'h1ff;
        mem[662] = 10'h3d3;
        mem[663] = 10'h394;
        mem[664] = 10'h33e;
        mem[665] = 10'h1a9;
        mem[666] = 10'h319;
        mem[667] = 10'h196;
        mem[668] = 10'h301;
        mem[669] = 10'h2e0;
        mem[670] = 10'h1e5;
        mem[671] = 10'h32c;
        mem[672] = 10'h0ed;
        mem[673] = 10'h36c;
        mem[674] = 10'h275;
        mem[675] = 10'h082;
        mem[676] = 10'h204;
        mem[677] = 10'h00c;
        mem[678] = 10'h1f4;
        mem[679] = 10'h3e3;
        mem[680] = 10'h1cd;
        mem[681] = 10'h38d;
        mem[682] = 10'h02b;
        mem[683] = 10'h257;
        mem[684] = 10'h18a;
        mem[685] = 10'h017;
        mem[686] = 10'h398;
        mem[687] = 10'h0ad;
        mem[688] = 10'h182;
        mem[689] = 10'h181;
        mem[690] = 10'h048;
        mem[691] = 10'h09a;
        mem[692] = 10'h3cf;
        mem[693] = 10'h294;
        mem[694] = 10'h2d4;
        mem[695] = 10'h1af;
        mem[696] = 10'h1b6;
        mem[697] = 10'h333;
        mem[698] = 10'h3d2;
        mem[699] = 10'h10a;
        mem[700] = 10'h28f;
        mem[701] = 10'h2c6;
        mem[702] = 10'h0ee;
        mem[703] = 10'h157;
        mem[704] = 10'h2f8;
        mem[705] = 10'h1db;
        mem[706] = 10'h079;
        mem[707] = 10'h3ab;
        mem[708] = 10'h2fc;
        mem[709] = 10'h0a1;
        mem[710] = 10'h1d8;
        mem[711] = 10'h27e;
        mem[712] = 10'h0cb;
        mem[713] = 10'h3c9;
        mem[714] = 10'h1b8;
        mem[715] = 10'h199;
        mem[716] = 10'h22a;
        mem[717] = 10'h358;
        mem[718] = 10'h328;
        mem[719] = 10'h3e8;
        mem[720] = 10'h326;
        mem[721] = 10'h058;
        mem[722] = 10'h12e;
        mem[723] = 10'h327;
        mem[724] = 10'h01d;
        mem[725] = 10'h3e4;
        mem[726] = 10'h26b;
        mem[727] = 10'h1a4;
        mem[728] = 10'h00d;
        mem[729] = 10'h33f;
        mem[730] = 10'h28a;
        mem[731] = 10'h32e;
        mem[732] = 10'h1b3;
        mem[733] = 10'h367;
        mem[734] = 10'h3cb;
        mem[735] = 10'h278;
        mem[736] = 10'h093;
        mem[737] = 10'h02a;
        mem[738] = 10'h3a6;
        mem[739] = 10'h0e7;
        mem[740] = 10'h02c;
        mem[741] = 10'h167;
        mem[742] = 10'h2c9;
        mem[743] = 10'h2ad;
        mem[744] = 10'h391;
        mem[745] = 10'h135;
        mem[746] = 10'h153;
        mem[747] = 10'h38e;
        mem[748] = 10'h36d;
        mem[749] = 10'h2a9;
        mem[750] = 10'h256;
        mem[751] = 10'h271;
        mem[752] = 10'h0a8;
        mem[753] = 10'h11a;
        mem[754] = 10'h2fb;
        mem[755] = 10'h3f2;
        mem[756] = 10'h096;
        mem[757] = 10'h0c1;
        mem[758] = 10'h389;
        mem[759] = 10'h109;
        mem[760] = 10'h3b8;
        mem[761] = 10'h1a6;
        mem[762] = 10'h2e5;
        mem[763] = 10'h304;
        mem[764] = 10'h055;
        mem[765] = 10'h0db;
        mem[766] = 10'h377;
        mem[767] = 10'h1ce;
        mem[768] = 10'h39b;
        mem[769] = 10'h13b;
        mem[770] = 10'h05f;
        mem[771] = 10'h05e;
        mem[772] = 10'h2ac;
        mem[773] = 10'h05d;
        mem[774] = 10'h074;
        mem[775] = 10'h280;
        mem[776] = 10'h3bb;
        mem[777] = 10'h325;
        mem[778] = 10'h07b;
        mem[779] = 10'h1fc;
        mem[780] = 10'h118;
        mem[781] = 10'h213;
        mem[782] = 10'h3d1;
        mem[783] = 10'h2d3;
        mem[784] = 10'h14d;
        mem[785] = 10'h174;
        mem[786] = 10'h0d6;
        mem[787] = 10'h121;
        mem[788] = 10'h08f;
        mem[789] = 10'h3b0;
        mem[790] = 10'h0f7;
        mem[791] = 10'h3da;
        mem[792] = 10'h0de;
        mem[793] = 10'h122;
        mem[794] = 10'h008;
        mem[795] = 10'h2b9;
        mem[796] = 10'h19d;
        mem[797] = 10'h3d4;
        mem[798] = 10'h3be;
        mem[799] = 10'h158;
        mem[800] = 10'h2c1;
        mem[801] = 10'h2f9;
        mem[802] = 10'h1ef;
        mem[803] = 10'h2bf;
        mem[804] = 10'h3ad;
        mem[805] = 10'h173;
        mem[806] = 10'h2a4;
        mem[807] = 10'h04c;
        mem[808] = 10'h138;
        mem[809] = 10'h3f0;
        mem[810] = 10'h1fb;
        mem[811] = 10'h151;
        mem[812] = 10'h2f1;
        mem[813] = 10'h0a2;
        mem[814] = 10'h286;
        mem[815] = 10'h075;
        mem[816] = 10'h3bf;
        mem[817] = 10'h3c8;
        mem[818] = 10'h08a;
        mem[819] = 10'h088;
        mem[820] = 10'h053;
        mem[821] = 10'h125;
        mem[822] = 10'h23a;
        mem[823] = 10'h07f;
        mem[824] = 10'h3df;
        mem[825] = 10'h038;
        mem[826] = 10'h384;
        mem[827] = 10'h0ce;
        mem[828] = 10'h165;
        mem[829] = 10'h019;
        mem[830] = 10'h312;
        mem[831] = 10'h139;
        mem[832] = 10'h24c;
        mem[833] = 10'h295;
        mem[834] = 10'h209;
        mem[835] = 10'h03a;
        mem[836] = 10'h1c1;
        mem[837] = 10'h317;
        mem[838] = 10'h2ff;
        mem[839] = 10'h13d;
        mem[840] = 10'h1bd;
        mem[841] = 10'h222;
        mem[842] = 10'h046;
        mem[843] = 10'h018;
        mem[844] = 10'h372;
        mem[845] = 10'h00b;
        mem[846] = 10'h34b;
        mem[847] = 10'h17b;
        mem[848] = 10'h20a;
        mem[849] = 10'h24a;
        mem[850] = 10'h3ed;
        mem[851] = 10'h22f;
        mem[852] = 10'h1d0;
        mem[853] = 10'h3b5;
        mem[854] = 10'h0bc;
        mem[855] = 10'h27d;
        mem[856] = 10'h06c;
        mem[857] = 10'h34c;
        mem[858] = 10'h087;
        mem[859] = 10'h11d;
        mem[860] = 10'h347;
        mem[861] = 10'h310;
        mem[862] = 10'h127;
        mem[863] = 10'h201;
        mem[864] = 10'h3eb;
        mem[865] = 10'h1b4;
        mem[866] = 10'h356;
        mem[867] = 10'h1bc;
        mem[868] = 10'h224;
        mem[869] = 10'h36b;
        mem[870] = 10'h064;
        mem[871] = 10'h355;
        mem[872] = 10'h0f8;
        mem[873] = 10'h290;
        mem[874] = 10'h1dc;
        mem[875] = 10'h129;
        mem[876] = 10'h080;
        mem[877] = 10'h236;
        mem[878] = 10'h1a5;
        mem[879] = 10'h2ea;
        mem[880] = 10'h1bb;
        mem[881] = 10'h251;
        mem[882] = 10'h2b3;
        mem[883] = 10'h1ec;
        mem[884] = 10'h175;
        mem[885] = 10'h133;
        mem[886] = 10'h35e;
        mem[887] = 10'h396;
        mem[888] = 10'h1fe;
        mem[889] = 10'h3a8;
        mem[890] = 10'h014;
        mem[891] = 10'h30f;
        mem[892] = 10'h24f;
        mem[893] = 10'h31e;
        mem[894] = 10'h1dd;
        mem[895] = 10'h1d2;
        mem[896] = 10'h02f;
        mem[897] = 10'h33d;
        mem[898] = 10'h2be;
        mem[899] = 10'h106;
        mem[900] = 10'h2f3;
        mem[901] = 10'h1ed;
        mem[902] = 10'h1e7;
        mem[903] = 10'h2cd;
        mem[904] = 10'h178;
        mem[905] = 10'h3bc;
        mem[906] = 10'h3b1;
        mem[907] = 10'h223;
        mem[908] = 10'h247;
        mem[909] = 10'h2e2;
        mem[910] = 10'h259;
        mem[911] = 10'h078;
        mem[912] = 10'h011;
        mem[913] = 10'h0b9;
        mem[914] = 10'h13f;
        mem[915] = 10'h244;
        mem[916] = 10'h09f;
        mem[917] = 10'h020;
        mem[918] = 10'h0c7;
        mem[919] = 10'h335;
        mem[920] = 10'h349;
        mem[921] = 10'h179;
        mem[922] = 10'h0e8;
        mem[923] = 10'h070;
        mem[924] = 10'h306;
        mem[925] = 10'h0c5;
        mem[926] = 10'h3fc;
        mem[927] = 10'h1b1;
        mem[928] = 10'h1c2;
        mem[929] = 10'h2f2;
        mem[930] = 10'h3ec;
        mem[931] = 10'h374;
        mem[932] = 10'h010;
        mem[933] = 10'h351;
        mem[934] = 10'h16b;
        mem[935] = 10'h28c;
        mem[936] = 10'h300;
        mem[937] = 10'h124;
        mem[938] = 10'h2f0;
        mem[939] = 10'h042;
        mem[940] = 10'h187;
        mem[941] = 10'h2b5;
        mem[942] = 10'h045;
        mem[943] = 10'h371;
        mem[944] = 10'h38c;
        mem[945] = 10'h2ce;
        mem[946] = 10'h06a;
        mem[947] = 10'h2ab;
        mem[948] = 10'h1f8;
        mem[949] = 10'h24d;
        mem[950] = 10'h2b7;
        mem[951] = 10'h253;
        mem[952] = 10'h1c0;
        mem[953] = 10'h3f4;
        mem[954] = 10'h321;
        mem[955] = 10'h0fd;
        mem[956] = 10'h0aa;
        mem[957] = 10'h094;
        mem[958] = 10'h193;
        mem[959] = 10'h051;
        mem[960] = 10'h0a0;
        mem[961] = 10'h21c;
        mem[962] = 10'h113;
        mem[963] = 10'h13e;
        mem[964] = 10'h375;
        mem[965] = 10'h08c;
        mem[966] = 10'h1a0;
        mem[967] = 10'h365;
        mem[968] = 10'h1d4;
        mem[969] = 10'h030;
        mem[970] = 10'h20d;
        mem[971] = 10'h363;
        mem[972] = 10'h237;
        mem[973] = 10'h0f4;
        mem[974] = 10'h318;
        mem[975] = 10'h026;
        mem[976] = 10'h3d5;
        mem[977] = 10'h104;
        mem[978] = 10'h188;
        mem[979] = 10'h14a;
        mem[980] = 10'h090;
        mem[981] = 10'h029;
        mem[982] = 10'h130;
        mem[983] = 10'h142;
        mem[984] = 10'h04e;
        mem[985] = 10'h231;
        mem[986] = 10'h31c;
        mem[987] = 10'h021;
        mem[988] = 10'h2b6;
        mem[989] = 10'h3b6;
        mem[990] = 10'h272;
        mem[991] = 10'h08e;
        mem[992] = 10'h07d;
        mem[993] = 10'h3c4;
        mem[994] = 10'h189;
        mem[995] = 10'h0d9;
        mem[996] = 10'h0b2;
        mem[997] = 10'h35f;
        mem[998] = 10'h098;
        mem[999] = 10'h381;
        mem[1000] = 10'h140;
        mem[1001] = 10'h159;
        mem[1002] = 10'h24b;
        mem[1003] = 10'h25d;
        mem[1004] = 10'h232;
        mem[1005] = 10'h2e8;
        mem[1006] = 10'h2fd;
        mem[1007] = 10'h245;
        mem[1008] = 10'h012;
        mem[1009] = 10'h35b;
        mem[1010] = 10'h32d;
        mem[1011] = 10'h11f;
        mem[1012] = 10'h1c3;
        mem[1013] = 10'h27a;
        mem[1014] = 10'h238;
        mem[1015] = 10'h378;
        mem[1016] = 10'h311;
        mem[1017] = 10'h17f;
        mem[1018] = 10'h0bb;
        mem[1019] = 10'h1ac;
        mem[1020] = 10'h2ed;
        mem[1021] = 10'h39d;
        mem[1022] = 10'h346;
        mem[1023] = 10'h3b4;
    end
endmodule

module odo_sbox_large7(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h1c2;
        mem[1] = 10'h133;
        mem[2] = 10'h009;
        mem[3] = 10'h230;
        mem[4] = 10'h33b;
        mem[5] = 10'h36b;
        mem[6] = 10'h0db;
        mem[7] = 10'h149;
        mem[8] = 10'h3f4;
        mem[9] = 10'h2b4;
        mem[10] = 10'h0c1;
        mem[11] = 10'h1ea;
        mem[12] = 10'h1d2;
        mem[13] = 10'h059;
        mem[14] = 10'h204;
        mem[15] = 10'h3c4;
        mem[16] = 10'h250;
        mem[17] = 10'h061;
        mem[18] = 10'h293;
        mem[19] = 10'h2db;
        mem[20] = 10'h277;
        mem[21] = 10'h333;
        mem[22] = 10'h0cd;
        mem[23] = 10'h083;
        mem[24] = 10'h0e8;
        mem[25] = 10'h2b9;
        mem[26] = 10'h143;
        mem[27] = 10'h242;
        mem[28] = 10'h36c;
        mem[29] = 10'h3e0;
        mem[30] = 10'h2ba;
        mem[31] = 10'h0e9;
        mem[32] = 10'h249;
        mem[33] = 10'h0b9;
        mem[34] = 10'h1dc;
        mem[35] = 10'h2a5;
        mem[36] = 10'h084;
        mem[37] = 10'h1c5;
        mem[38] = 10'h259;
        mem[39] = 10'h2f2;
        mem[40] = 10'h38b;
        mem[41] = 10'h174;
        mem[42] = 10'h304;
        mem[43] = 10'h1f4;
        mem[44] = 10'h0cc;
        mem[45] = 10'h068;
        mem[46] = 10'h27b;
        mem[47] = 10'h3f1;
        mem[48] = 10'h3a1;
        mem[49] = 10'h186;
        mem[50] = 10'h380;
        mem[51] = 10'h1e7;
        mem[52] = 10'h229;
        mem[53] = 10'h311;
        mem[54] = 10'h0d0;
        mem[55] = 10'h1fe;
        mem[56] = 10'h134;
        mem[57] = 10'h0a6;
        mem[58] = 10'h2da;
        mem[59] = 10'h02d;
        mem[60] = 10'h001;
        mem[61] = 10'h3d6;
        mem[62] = 10'h37f;
        mem[63] = 10'h18a;
        mem[64] = 10'h065;
        mem[65] = 10'h15c;
        mem[66] = 10'h240;
        mem[67] = 10'h071;
        mem[68] = 10'h05b;
        mem[69] = 10'h02c;
        mem[70] = 10'h21f;
        mem[71] = 10'h090;
        mem[72] = 10'h39c;
        mem[73] = 10'h10b;
        mem[74] = 10'h3c1;
        mem[75] = 10'h334;
        mem[76] = 10'h1f7;
        mem[77] = 10'h0ac;
        mem[78] = 10'h1a9;
        mem[79] = 10'h1e2;
        mem[80] = 10'h02e;
        mem[81] = 10'h119;
        mem[82] = 10'h31c;
        mem[83] = 10'h2a1;
        mem[84] = 10'h3b4;
        mem[85] = 10'h2bf;
        mem[86] = 10'h371;
        mem[87] = 10'h087;
        mem[88] = 10'h00b;
        mem[89] = 10'h346;
        mem[90] = 10'h142;
        mem[91] = 10'h2d0;
        mem[92] = 10'h166;
        mem[93] = 10'h0bd;
        mem[94] = 10'h012;
        mem[95] = 10'h03a;
        mem[96] = 10'h226;
        mem[97] = 10'h2d2;
        mem[98] = 10'h393;
        mem[99] = 10'h2d7;
        mem[100] = 10'h38c;
        mem[101] = 10'h15f;
        mem[102] = 10'h081;
        mem[103] = 10'h01c;
        mem[104] = 10'h00e;
        mem[105] = 10'h2b5;
        mem[106] = 10'h252;
        mem[107] = 10'h348;
        mem[108] = 10'h121;
        mem[109] = 10'h2d4;
        mem[110] = 10'h197;
        mem[111] = 10'h07b;
        mem[112] = 10'h109;
        mem[113] = 10'h0f1;
        mem[114] = 10'h01a;
        mem[115] = 10'h247;
        mem[116] = 10'h2d8;
        mem[117] = 10'h3d9;
        mem[118] = 10'h20b;
        mem[119] = 10'h06b;
        mem[120] = 10'h0a7;
        mem[121] = 10'h18c;
        mem[122] = 10'h0d8;
        mem[123] = 10'h2ae;
        mem[124] = 10'h35c;
        mem[125] = 10'h152;
        mem[126] = 10'h215;
        mem[127] = 10'h363;
        mem[128] = 10'h32b;
        mem[129] = 10'h322;
        mem[130] = 10'h1ee;
        mem[131] = 10'h1ba;
        mem[132] = 10'h12c;
        mem[133] = 10'h1c1;
        mem[134] = 10'h206;
        mem[135] = 10'h01f;
        mem[136] = 10'h21c;
        mem[137] = 10'h236;
        mem[138] = 10'h0c5;
        mem[139] = 10'h23e;
        mem[140] = 10'h2e0;
        mem[141] = 10'h28b;
        mem[142] = 10'h3ec;
        mem[143] = 10'h22c;
        mem[144] = 10'h3ea;
        mem[145] = 10'h3ac;
        mem[146] = 10'h369;
        mem[147] = 10'h31a;
        mem[148] = 10'h060;
        mem[149] = 10'h307;
        mem[150] = 10'h26d;
        mem[151] = 10'h251;
        mem[152] = 10'h086;
        mem[153] = 10'h235;
        mem[154] = 10'h2f7;
        mem[155] = 10'h013;
        mem[156] = 10'h37a;
        mem[157] = 10'h38a;
        mem[158] = 10'h17b;
        mem[159] = 10'h13e;
        mem[160] = 10'h3bd;
        mem[161] = 10'h2d5;
        mem[162] = 10'h395;
        mem[163] = 10'h0f8;
        mem[164] = 10'h22d;
        mem[165] = 10'h002;
        mem[166] = 10'h3fd;
        mem[167] = 10'h256;
        mem[168] = 10'h248;
        mem[169] = 10'h201;
        mem[170] = 10'h0d7;
        mem[171] = 10'h35f;
        mem[172] = 10'h22e;
        mem[173] = 10'h366;
        mem[174] = 10'h20c;
        mem[175] = 10'h1eb;
        mem[176] = 10'h3e9;
        mem[177] = 10'h253;
        mem[178] = 10'h298;
        mem[179] = 10'h3bc;
        mem[180] = 10'h097;
        mem[181] = 10'h3a6;
        mem[182] = 10'h31d;
        mem[183] = 10'h397;
        mem[184] = 10'h0ce;
        mem[185] = 10'h138;
        mem[186] = 10'h23f;
        mem[187] = 10'h0fa;
        mem[188] = 10'h282;
        mem[189] = 10'h29a;
        mem[190] = 10'h1de;
        mem[191] = 10'h1d4;
        mem[192] = 10'h1da;
        mem[193] = 10'h241;
        mem[194] = 10'h3db;
        mem[195] = 10'h1ae;
        mem[196] = 10'h16e;
        mem[197] = 10'h3ff;
        mem[198] = 10'h1e8;
        mem[199] = 10'h2dc;
        mem[200] = 10'h191;
        mem[201] = 10'h302;
        mem[202] = 10'h356;
        mem[203] = 10'h06c;
        mem[204] = 10'h1a6;
        mem[205] = 10'h2ea;
        mem[206] = 10'h244;
        mem[207] = 10'h385;
        mem[208] = 10'h127;
        mem[209] = 10'h177;
        mem[210] = 10'h0fc;
        mem[211] = 10'h0c3;
        mem[212] = 10'h228;
        mem[213] = 10'h3ce;
        mem[214] = 10'h106;
        mem[215] = 10'h05f;
        mem[216] = 10'h11d;
        mem[217] = 10'h2e2;
        mem[218] = 10'h233;
        mem[219] = 10'h05c;
        mem[220] = 10'h3cb;
        mem[221] = 10'h3cf;
        mem[222] = 10'h18e;
        mem[223] = 10'h20e;
        mem[224] = 10'h056;
        mem[225] = 10'h118;
        mem[226] = 10'h100;
        mem[227] = 10'h113;
        mem[228] = 10'h0ef;
        mem[229] = 10'h0b4;
        mem[230] = 10'h0b5;
        mem[231] = 10'h224;
        mem[232] = 10'h155;
        mem[233] = 10'h1b8;
        mem[234] = 10'h089;
        mem[235] = 10'h1d8;
        mem[236] = 10'h26e;
        mem[237] = 10'h095;
        mem[238] = 10'h15d;
        mem[239] = 10'h299;
        mem[240] = 10'h123;
        mem[241] = 10'h159;
        mem[242] = 10'h1af;
        mem[243] = 10'h2a7;
        mem[244] = 10'h04a;
        mem[245] = 10'h09f;
        mem[246] = 10'h183;
        mem[247] = 10'h189;
        mem[248] = 10'h077;
        mem[249] = 10'h0e7;
        mem[250] = 10'h2f0;
        mem[251] = 10'h050;
        mem[252] = 10'h1d6;
        mem[253] = 10'h00c;
        mem[254] = 10'h368;
        mem[255] = 10'h303;
        mem[256] = 10'h29e;
        mem[257] = 10'h1be;
        mem[258] = 10'h386;
        mem[259] = 10'h00a;
        mem[260] = 10'h0c8;
        mem[261] = 10'h2c7;
        mem[262] = 10'h196;
        mem[263] = 10'h3f9;
        mem[264] = 10'h173;
        mem[265] = 10'h066;
        mem[266] = 10'h1dd;
        mem[267] = 10'h161;
        mem[268] = 10'h044;
        mem[269] = 10'h015;
        mem[270] = 10'h04c;
        mem[271] = 10'h0df;
        mem[272] = 10'h266;
        mem[273] = 10'h257;
        mem[274] = 10'h2b8;
        mem[275] = 10'h2e8;
        mem[276] = 10'h246;
        mem[277] = 10'h3b0;
        mem[278] = 10'h378;
        mem[279] = 10'h03c;
        mem[280] = 10'h0de;
        mem[281] = 10'h1f5;
        mem[282] = 10'h23d;
        mem[283] = 10'h17d;
        mem[284] = 10'h129;
        mem[285] = 10'h1df;
        mem[286] = 10'h23c;
        mem[287] = 10'h1f8;
        mem[288] = 10'h36d;
        mem[289] = 10'h376;
        mem[290] = 10'h192;
        mem[291] = 10'h31b;
        mem[292] = 10'h1ed;
        mem[293] = 10'h283;
        mem[294] = 10'h278;
        mem[295] = 10'h04d;
        mem[296] = 10'h007;
        mem[297] = 10'h157;
        mem[298] = 10'h1b9;
        mem[299] = 10'h067;
        mem[300] = 10'h0f6;
        mem[301] = 10'h2c0;
        mem[302] = 10'h1fd;
        mem[303] = 10'h026;
        mem[304] = 10'h14b;
        mem[305] = 10'h3c0;
        mem[306] = 10'h1e6;
        mem[307] = 10'h0c0;
        mem[308] = 10'h0fb;
        mem[309] = 10'h273;
        mem[310] = 10'h19b;
        mem[311] = 10'h19f;
        mem[312] = 10'h008;
        mem[313] = 10'h130;
        mem[314] = 10'h222;
        mem[315] = 10'h0e6;
        mem[316] = 10'h005;
        mem[317] = 10'h28c;
        mem[318] = 10'h13d;
        mem[319] = 10'h1c4;
        mem[320] = 10'h075;
        mem[321] = 10'h031;
        mem[322] = 10'h076;
        mem[323] = 10'h0b7;
        mem[324] = 10'h313;
        mem[325] = 10'h1bb;
        mem[326] = 10'h25d;
        mem[327] = 10'h1c7;
        mem[328] = 10'h0a5;
        mem[329] = 10'h010;
        mem[330] = 10'h312;
        mem[331] = 10'h284;
        mem[332] = 10'h0bf;
        mem[333] = 10'h073;
        mem[334] = 10'h29d;
        mem[335] = 10'h382;
        mem[336] = 10'h0e3;
        mem[337] = 10'h1d9;
        mem[338] = 10'h1e0;
        mem[339] = 10'h1e3;
        mem[340] = 10'h1ff;
        mem[341] = 10'h30e;
        mem[342] = 10'h287;
        mem[343] = 10'h340;
        mem[344] = 10'h1d3;
        mem[345] = 10'h025;
        mem[346] = 10'h3a7;
        mem[347] = 10'h25a;
        mem[348] = 10'h32f;
        mem[349] = 10'h12e;
        mem[350] = 10'h383;
        mem[351] = 10'h037;
        mem[352] = 10'h28e;
        mem[353] = 10'h0d4;
        mem[354] = 10'h315;
        mem[355] = 10'h2f3;
        mem[356] = 10'h2c5;
        mem[357] = 10'h35a;
        mem[358] = 10'h1d5;
        mem[359] = 10'h3b1;
        mem[360] = 10'h07c;
        mem[361] = 10'h1cd;
        mem[362] = 10'h1c0;
        mem[363] = 10'h2ee;
        mem[364] = 10'h306;
        mem[365] = 10'h34d;
        mem[366] = 10'h342;
        mem[367] = 10'h3f8;
        mem[368] = 10'h111;
        mem[369] = 10'h3ee;
        mem[370] = 10'h29c;
        mem[371] = 10'h1a2;
        mem[372] = 10'h210;
        mem[373] = 10'h211;
        mem[374] = 10'h3ae;
        mem[375] = 10'h171;
        mem[376] = 10'h2c6;
        mem[377] = 10'h338;
        mem[378] = 10'h26f;
        mem[379] = 10'h238;
        mem[380] = 10'h361;
        mem[381] = 10'h1fa;
        mem[382] = 10'h064;
        mem[383] = 10'h09c;
        mem[384] = 10'h219;
        mem[385] = 10'h2cb;
        mem[386] = 10'h349;
        mem[387] = 10'h2cf;
        mem[388] = 10'h243;
        mem[389] = 10'h058;
        mem[390] = 10'h132;
        mem[391] = 10'h245;
        mem[392] = 10'h30b;
        mem[393] = 10'h22a;
        mem[394] = 10'h30f;
        mem[395] = 10'h09d;
        mem[396] = 10'h2b3;
        mem[397] = 10'h131;
        mem[398] = 10'h05d;
        mem[399] = 10'h21e;
        mem[400] = 10'h179;
        mem[401] = 10'h263;
        mem[402] = 10'h17e;
        mem[403] = 10'h027;
        mem[404] = 10'h020;
        mem[405] = 10'h1f6;
        mem[406] = 10'h212;
        mem[407] = 10'h190;
        mem[408] = 10'h300;
        mem[409] = 10'h202;
        mem[410] = 10'h114;
        mem[411] = 10'h35d;
        mem[412] = 10'h364;
        mem[413] = 10'h162;
        mem[414] = 10'h267;
        mem[415] = 10'h006;
        mem[416] = 10'h32e;
        mem[417] = 10'h3aa;
        mem[418] = 10'h362;
        mem[419] = 10'h38f;
        mem[420] = 10'h0a4;
        mem[421] = 10'h0be;
        mem[422] = 10'h272;
        mem[423] = 10'h0b8;
        mem[424] = 10'h24e;
        mem[425] = 10'h1a4;
        mem[426] = 10'h115;
        mem[427] = 10'h3c2;
        mem[428] = 10'h1db;
        mem[429] = 10'h137;
        mem[430] = 10'h0a1;
        mem[431] = 10'h2ac;
        mem[432] = 10'h33c;
        mem[433] = 10'h264;
        mem[434] = 10'h3a9;
        mem[435] = 10'h035;
        mem[436] = 10'h254;
        mem[437] = 10'h03e;
        mem[438] = 10'h1fc;
        mem[439] = 10'h22f;
        mem[440] = 10'h107;
        mem[441] = 10'h003;
        mem[442] = 10'h331;
        mem[443] = 10'h182;
        mem[444] = 10'h181;
        mem[445] = 10'h261;
        mem[446] = 10'h135;
        mem[447] = 10'h345;
        mem[448] = 10'h3fe;
        mem[449] = 10'h387;
        mem[450] = 10'h375;
        mem[451] = 10'h12d;
        mem[452] = 10'h37c;
        mem[453] = 10'h185;
        mem[454] = 10'h317;
        mem[455] = 10'h2d1;
        mem[456] = 10'h018;
        mem[457] = 10'h11a;
        mem[458] = 10'h39a;
        mem[459] = 10'h3d0;
        mem[460] = 10'h102;
        mem[461] = 10'h351;
        mem[462] = 10'h398;
        mem[463] = 10'h085;
        mem[464] = 10'h0dc;
        mem[465] = 10'h3cd;
        mem[466] = 10'h2ab;
        mem[467] = 10'h0d9;
        mem[468] = 10'h269;
        mem[469] = 10'h0f4;
        mem[470] = 10'h285;
        mem[471] = 10'h1b7;
        mem[472] = 10'h2a9;
        mem[473] = 10'h3b8;
        mem[474] = 10'h357;
        mem[475] = 10'h27e;
        mem[476] = 10'h0eb;
        mem[477] = 10'h36f;
        mem[478] = 10'h2ef;
        mem[479] = 10'h2a6;
        mem[480] = 10'h10e;
        mem[481] = 10'h341;
        mem[482] = 10'h255;
        mem[483] = 10'h3de;
        mem[484] = 10'h12f;
        mem[485] = 10'h1cb;
        mem[486] = 10'h1b2;
        mem[487] = 10'h24f;
        mem[488] = 10'h1a0;
        mem[489] = 10'h033;
        mem[490] = 10'h180;
        mem[491] = 10'h21a;
        mem[492] = 10'h2af;
        mem[493] = 10'h27d;
        mem[494] = 10'h0ae;
        mem[495] = 10'h326;
        mem[496] = 10'h0a3;
        mem[497] = 10'h3d3;
        mem[498] = 10'h124;
        mem[499] = 10'h0b3;
        mem[500] = 10'h268;
        mem[501] = 10'h39b;
        mem[502] = 10'h07a;
        mem[503] = 10'h04b;
        mem[504] = 10'h04f;
        mem[505] = 10'h3e6;
        mem[506] = 10'h328;
        mem[507] = 10'h3e5;
        mem[508] = 10'h354;
        mem[509] = 10'h19e;
        mem[510] = 10'h110;
        mem[511] = 10'h141;
        mem[512] = 10'h163;
        mem[513] = 10'h101;
        mem[514] = 10'h344;
        mem[515] = 10'h0fd;
        mem[516] = 10'h0a0;
        mem[517] = 10'h049;
        mem[518] = 10'h108;
        mem[519] = 10'h1a7;
        mem[520] = 10'h3d5;
        mem[521] = 10'h3bf;
        mem[522] = 10'h360;
        mem[523] = 10'h205;
        mem[524] = 10'h365;
        mem[525] = 10'h26b;
        mem[526] = 10'h21b;
        mem[527] = 10'h1ef;
        mem[528] = 10'h225;
        mem[529] = 10'h2b0;
        mem[530] = 10'h08d;
        mem[531] = 10'h271;
        mem[532] = 10'h004;
        mem[533] = 10'h116;
        mem[534] = 10'h27c;
        mem[535] = 10'h231;
        mem[536] = 10'h3a5;
        mem[537] = 10'h0b2;
        mem[538] = 10'h379;
        mem[539] = 10'h0a8;
        mem[540] = 10'h1c8;
        mem[541] = 10'h3f3;
        mem[542] = 10'h06f;
        mem[543] = 10'h1c6;
        mem[544] = 10'h136;
        mem[545] = 10'h045;
        mem[546] = 10'h08b;
        mem[547] = 10'h14a;
        mem[548] = 10'h1c3;
        mem[549] = 10'h2c2;
        mem[550] = 10'h1b0;
        mem[551] = 10'h3ab;
        mem[552] = 10'h20a;
        mem[553] = 10'h24c;
        mem[554] = 10'h11e;
        mem[555] = 10'h151;
        mem[556] = 10'h1a5;
        mem[557] = 10'h3dd;
        mem[558] = 10'h2fc;
        mem[559] = 10'h17a;
        mem[560] = 10'h394;
        mem[561] = 10'h09e;
        mem[562] = 10'h0cf;
        mem[563] = 10'h276;
        mem[564] = 10'h0aa;
        mem[565] = 10'h358;
        mem[566] = 10'h150;
        mem[567] = 10'h25b;
        mem[568] = 10'h2e3;
        mem[569] = 10'h147;
        mem[570] = 10'h234;
        mem[571] = 10'h092;
        mem[572] = 10'h082;
        mem[573] = 10'h07d;
        mem[574] = 10'h3e4;
        mem[575] = 10'h0c9;
        mem[576] = 10'h11f;
        mem[577] = 10'h0ba;
        mem[578] = 10'h0ed;
        mem[579] = 10'h2d9;
        mem[580] = 10'h10f;
        mem[581] = 10'h088;
        mem[582] = 10'h169;
        mem[583] = 10'h0d3;
        mem[584] = 10'h3cc;
        mem[585] = 10'h03d;
        mem[586] = 10'h04e;
        mem[587] = 10'h09b;
        mem[588] = 10'h2fa;
        mem[589] = 10'h319;
        mem[590] = 10'h2e5;
        mem[591] = 10'h1e5;
        mem[592] = 10'h34e;
        mem[593] = 10'h2fd;
        mem[594] = 10'h14d;
        mem[595] = 10'h0a2;
        mem[596] = 10'h14c;
        mem[597] = 10'h213;
        mem[598] = 10'h024;
        mem[599] = 10'h0cb;
        mem[600] = 10'h33e;
        mem[601] = 10'h093;
        mem[602] = 10'h15b;
        mem[603] = 10'h06d;
        mem[604] = 10'h3da;
        mem[605] = 10'h314;
        mem[606] = 10'h062;
        mem[607] = 10'h167;
        mem[608] = 10'h2d3;
        mem[609] = 10'h23b;
        mem[610] = 10'h396;
        mem[611] = 10'h31f;
        mem[612] = 10'h34b;
        mem[613] = 10'h139;
        mem[614] = 10'h3c6;
        mem[615] = 10'h08f;
        mem[616] = 10'h18b;
        mem[617] = 10'h28a;
        mem[618] = 10'h329;
        mem[619] = 10'h1c9;
        mem[620] = 10'h16a;
        mem[621] = 10'h0b6;
        mem[622] = 10'h098;
        mem[623] = 10'h16b;
        mem[624] = 10'h399;
        mem[625] = 10'h353;
        mem[626] = 10'h218;
        mem[627] = 10'h188;
        mem[628] = 10'h3fc;
        mem[629] = 10'h0e4;
        mem[630] = 10'h126;
        mem[631] = 10'h3be;
        mem[632] = 10'h2b1;
        mem[633] = 10'h0f0;
        mem[634] = 10'h014;
        mem[635] = 10'h01d;
        mem[636] = 10'h0e2;
        mem[637] = 10'h184;
        mem[638] = 10'h023;
        mem[639] = 10'h2ca;
        mem[640] = 10'h156;
        mem[641] = 10'h28f;
        mem[642] = 10'h3a0;
        mem[643] = 10'h3a3;
        mem[644] = 10'h1f1;
        mem[645] = 10'h24a;
        mem[646] = 10'h022;
        mem[647] = 10'h37e;
        mem[648] = 10'h13b;
        mem[649] = 10'h2e6;
        mem[650] = 10'h296;
        mem[651] = 10'h145;
        mem[652] = 10'h223;
        mem[653] = 10'h178;
        mem[654] = 10'h096;
        mem[655] = 10'h122;
        mem[656] = 10'h07e;
        mem[657] = 10'h029;
        mem[658] = 10'h24d;
        mem[659] = 10'h3ef;
        mem[660] = 10'h3f5;
        mem[661] = 10'h2cd;
        mem[662] = 10'h10a;
        mem[663] = 10'h347;
        mem[664] = 10'h2a0;
        mem[665] = 10'h289;
        mem[666] = 10'h3dc;
        mem[667] = 10'h200;
        mem[668] = 10'h37d;
        mem[669] = 10'h2fe;
        mem[670] = 10'h0d6;
        mem[671] = 10'h3a2;
        mem[672] = 10'h232;
        mem[673] = 10'h154;
        mem[674] = 10'h335;
        mem[675] = 10'h208;
        mem[676] = 10'h07f;
        mem[677] = 10'h18d;
        mem[678] = 10'h3b3;
        mem[679] = 10'h1b4;
        mem[680] = 10'h330;
        mem[681] = 10'h000;
        mem[682] = 10'h281;
        mem[683] = 10'h0d1;
        mem[684] = 10'h270;
        mem[685] = 10'h275;
        mem[686] = 10'h209;
        mem[687] = 10'h06a;
        mem[688] = 10'h26c;
        mem[689] = 10'h1bd;
        mem[690] = 10'h3b6;
        mem[691] = 10'h0b0;
        mem[692] = 10'h0ec;
        mem[693] = 10'h2b7;
        mem[694] = 10'h038;
        mem[695] = 10'h105;
        mem[696] = 10'h12b;
        mem[697] = 10'h350;
        mem[698] = 10'h1e1;
        mem[699] = 10'h1a1;
        mem[700] = 10'h195;
        mem[701] = 10'h13f;
        mem[702] = 10'h078;
        mem[703] = 10'h3d4;
        mem[704] = 10'h1ce;
        mem[705] = 10'h055;
        mem[706] = 10'h2f9;
        mem[707] = 10'h3d7;
        mem[708] = 10'h16f;
        mem[709] = 10'h0f3;
        mem[710] = 10'h2ec;
        mem[711] = 10'h2e1;
        mem[712] = 10'h390;
        mem[713] = 10'h041;
        mem[714] = 10'h217;
        mem[715] = 10'h0ff;
        mem[716] = 10'h165;
        mem[717] = 10'h3a8;
        mem[718] = 10'h144;
        mem[719] = 10'h0c6;
        mem[720] = 10'h016;
        mem[721] = 10'h01e;
        mem[722] = 10'h332;
        mem[723] = 10'h3b5;
        mem[724] = 10'h1bc;
        mem[725] = 10'h343;
        mem[726] = 10'h3d1;
        mem[727] = 10'h216;
        mem[728] = 10'h15a;
        mem[729] = 10'h260;
        mem[730] = 10'h3ca;
        mem[731] = 10'h2f5;
        mem[732] = 10'h33a;
        mem[733] = 10'h31e;
        mem[734] = 10'h0c2;
        mem[735] = 10'h13a;
        mem[736] = 10'h32c;
        mem[737] = 10'h08a;
        mem[738] = 10'h38d;
        mem[739] = 10'h0bc;
        mem[740] = 10'h12a;
        mem[741] = 10'h0af;
        mem[742] = 10'h279;
        mem[743] = 10'h3ed;
        mem[744] = 10'h392;
        mem[745] = 10'h14f;
        mem[746] = 10'h094;
        mem[747] = 10'h3b7;
        mem[748] = 10'h2be;
        mem[749] = 10'h046;
        mem[750] = 10'h172;
        mem[751] = 10'h310;
        mem[752] = 10'h2dd;
        mem[753] = 10'h176;
        mem[754] = 10'h262;
        mem[755] = 10'h148;
        mem[756] = 10'h374;
        mem[757] = 10'h2c9;
        mem[758] = 10'h2f8;
        mem[759] = 10'h372;
        mem[760] = 10'h048;
        mem[761] = 10'h29f;
        mem[762] = 10'h19d;
        mem[763] = 10'h227;
        mem[764] = 10'h3f2;
        mem[765] = 10'h0ea;
        mem[766] = 10'h3e2;
        mem[767] = 10'h05e;
        mem[768] = 10'h074;
        mem[769] = 10'h258;
        mem[770] = 10'h02b;
        mem[771] = 10'h128;
        mem[772] = 10'h070;
        mem[773] = 10'h2e4;
        mem[774] = 10'h0e0;
        mem[775] = 10'h0f9;
        mem[776] = 10'h336;
        mem[777] = 10'h23a;
        mem[778] = 10'h1bf;
        mem[779] = 10'h355;
        mem[780] = 10'h27a;
        mem[781] = 10'h16d;
        mem[782] = 10'h3af;
        mem[783] = 10'h198;
        mem[784] = 10'h099;
        mem[785] = 10'h1b6;
        mem[786] = 10'h2ed;
        mem[787] = 10'h288;
        mem[788] = 10'h0d5;
        mem[789] = 10'h112;
        mem[790] = 10'h34f;
        mem[791] = 10'h2a8;
        mem[792] = 10'h1f2;
        mem[793] = 10'h34a;
        mem[794] = 10'h3b2;
        mem[795] = 10'h011;
        mem[796] = 10'h01b;
        mem[797] = 10'h39d;
        mem[798] = 10'h1d1;
        mem[799] = 10'h22b;
        mem[800] = 10'h3bb;
        mem[801] = 10'h2c4;
        mem[802] = 10'h35e;
        mem[803] = 10'h187;
        mem[804] = 10'h054;
        mem[805] = 10'h318;
        mem[806] = 10'h1fb;
        mem[807] = 10'h052;
        mem[808] = 10'h30d;
        mem[809] = 10'h03f;
        mem[810] = 10'h09a;
        mem[811] = 10'h26a;
        mem[812] = 10'h21d;
        mem[813] = 10'h039;
        mem[814] = 10'h1d0;
        mem[815] = 10'h1f0;
        mem[816] = 10'h34c;
        mem[817] = 10'h028;
        mem[818] = 10'h3c7;
        mem[819] = 10'h295;
        mem[820] = 10'h36e;
        mem[821] = 10'h207;
        mem[822] = 10'h38e;
        mem[823] = 10'h091;
        mem[824] = 10'h3f0;
        mem[825] = 10'h377;
        mem[826] = 10'h199;
        mem[827] = 10'h117;
        mem[828] = 10'h158;
        mem[829] = 10'h2de;
        mem[830] = 10'h25e;
        mem[831] = 10'h3a4;
        mem[832] = 10'h384;
        mem[833] = 10'h11c;
        mem[834] = 10'h168;
        mem[835] = 10'h239;
        mem[836] = 10'h20d;
        mem[837] = 10'h2aa;
        mem[838] = 10'h1f9;
        mem[839] = 10'h265;
        mem[840] = 10'h373;
        mem[841] = 10'h2d6;
        mem[842] = 10'h3c5;
        mem[843] = 10'h08e;
        mem[844] = 10'h3df;
        mem[845] = 10'h1b5;
        mem[846] = 10'h286;
        mem[847] = 10'h29b;
        mem[848] = 10'h25c;
        mem[849] = 10'h2b2;
        mem[850] = 10'h28d;
        mem[851] = 10'h290;
        mem[852] = 10'h3f7;
        mem[853] = 10'h160;
        mem[854] = 10'h3e3;
        mem[855] = 10'h2b6;
        mem[856] = 10'h034;
        mem[857] = 10'h040;
        mem[858] = 10'h2f4;
        mem[859] = 10'h15e;
        mem[860] = 10'h3c3;
        mem[861] = 10'h16c;
        mem[862] = 10'h370;
        mem[863] = 10'h1a3;
        mem[864] = 10'h2bc;
        mem[865] = 10'h0f5;
        mem[866] = 10'h291;
        mem[867] = 10'h0d2;
        mem[868] = 10'h0fe;
        mem[869] = 10'h3ba;
        mem[870] = 10'h19a;
        mem[871] = 10'h274;
        mem[872] = 10'h20f;
        mem[873] = 10'h2f6;
        mem[874] = 10'h3e7;
        mem[875] = 10'h063;
        mem[876] = 10'h391;
        mem[877] = 10'h069;
        mem[878] = 10'h02f;
        mem[879] = 10'h1ca;
        mem[880] = 10'h3fb;
        mem[881] = 10'h325;
        mem[882] = 10'h2ff;
        mem[883] = 10'h0ad;
        mem[884] = 10'h019;
        mem[885] = 10'h194;
        mem[886] = 10'h14e;
        mem[887] = 10'h327;
        mem[888] = 10'h367;
        mem[889] = 10'h359;
        mem[890] = 10'h021;
        mem[891] = 10'h2f1;
        mem[892] = 10'h1e4;
        mem[893] = 10'h1cc;
        mem[894] = 10'h280;
        mem[895] = 10'h1ad;
        mem[896] = 10'h1e9;
        mem[897] = 10'h37b;
        mem[898] = 10'h053;
        mem[899] = 10'h3e8;
        mem[900] = 10'h1ec;
        mem[901] = 10'h072;
        mem[902] = 10'h292;
        mem[903] = 10'h1ab;
        mem[904] = 10'h125;
        mem[905] = 10'h00f;
        mem[906] = 10'h104;
        mem[907] = 10'h2eb;
        mem[908] = 10'h140;
        mem[909] = 10'h221;
        mem[910] = 10'h2e9;
        mem[911] = 10'h1aa;
        mem[912] = 10'h043;
        mem[913] = 10'h3fa;
        mem[914] = 10'h25f;
        mem[915] = 10'h103;
        mem[916] = 10'h0ab;
        mem[917] = 10'h39f;
        mem[918] = 10'h3c8;
        mem[919] = 10'h2a2;
        mem[920] = 10'h120;
        mem[921] = 10'h03b;
        mem[922] = 10'h10c;
        mem[923] = 10'h17f;
        mem[924] = 10'h1b1;
        mem[925] = 10'h0ee;
        mem[926] = 10'h1d7;
        mem[927] = 10'h1f3;
        mem[928] = 10'h3f6;
        mem[929] = 10'h193;
        mem[930] = 10'h00d;
        mem[931] = 10'h047;
        mem[932] = 10'h2a3;
        mem[933] = 10'h042;
        mem[934] = 10'h2a4;
        mem[935] = 10'h17c;
        mem[936] = 10'h08c;
        mem[937] = 10'h079;
        mem[938] = 10'h017;
        mem[939] = 10'h339;
        mem[940] = 10'h0f7;
        mem[941] = 10'h1cf;
        mem[942] = 10'h320;
        mem[943] = 10'h3e1;
        mem[944] = 10'h19c;
        mem[945] = 10'h27f;
        mem[946] = 10'h337;
        mem[947] = 10'h032;
        mem[948] = 10'h294;
        mem[949] = 10'h080;
        mem[950] = 10'h0dd;
        mem[951] = 10'h10d;
        mem[952] = 10'h297;
        mem[953] = 10'h2cc;
        mem[954] = 10'h02a;
        mem[955] = 10'h24b;
        mem[956] = 10'h30c;
        mem[957] = 10'h324;
        mem[958] = 10'h2bd;
        mem[959] = 10'h13c;
        mem[960] = 10'h0b1;
        mem[961] = 10'h11b;
        mem[962] = 10'h220;
        mem[963] = 10'h237;
        mem[964] = 10'h35b;
        mem[965] = 10'h2fb;
        mem[966] = 10'h301;
        mem[967] = 10'h323;
        mem[968] = 10'h2ad;
        mem[969] = 10'h3d2;
        mem[970] = 10'h0e1;
        mem[971] = 10'h2df;
        mem[972] = 10'h2c3;
        mem[973] = 10'h05a;
        mem[974] = 10'h030;
        mem[975] = 10'h309;
        mem[976] = 10'h1ac;
        mem[977] = 10'h2c8;
        mem[978] = 10'h3d8;
        mem[979] = 10'h308;
        mem[980] = 10'h1b3;
        mem[981] = 10'h2c1;
        mem[982] = 10'h146;
        mem[983] = 10'h32a;
        mem[984] = 10'h3b9;
        mem[985] = 10'h203;
        mem[986] = 10'h352;
        mem[987] = 10'h2bb;
        mem[988] = 10'h388;
        mem[989] = 10'h0ca;
        mem[990] = 10'h316;
        mem[991] = 10'h2ce;
        mem[992] = 10'h39e;
        mem[993] = 10'h3eb;
        mem[994] = 10'h36a;
        mem[995] = 10'h0a9;
        mem[996] = 10'h057;
        mem[997] = 10'h0e5;
        mem[998] = 10'h305;
        mem[999] = 10'h0da;
        mem[1000] = 10'h214;
        mem[1001] = 10'h18f;
        mem[1002] = 10'h2e7;
        mem[1003] = 10'h06e;
        mem[1004] = 10'h30a;
        mem[1005] = 10'h051;
        mem[1006] = 10'h1a8;
        mem[1007] = 10'h3c9;
        mem[1008] = 10'h0bb;
        mem[1009] = 10'h389;
        mem[1010] = 10'h33d;
        mem[1011] = 10'h175;
        mem[1012] = 10'h381;
        mem[1013] = 10'h036;
        mem[1014] = 10'h33f;
        mem[1015] = 10'h164;
        mem[1016] = 10'h170;
        mem[1017] = 10'h3ad;
        mem[1018] = 10'h153;
        mem[1019] = 10'h32d;
        mem[1020] = 10'h321;
        mem[1021] = 10'h0c4;
        mem[1022] = 10'h0c7;
        mem[1023] = 10'h0f2;
    end
endmodule

module odo_sbox_large8(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h207;
        mem[1] = 10'h38b;
        mem[2] = 10'h3fd;
        mem[3] = 10'h2fe;
        mem[4] = 10'h36f;
        mem[5] = 10'h0f8;
        mem[6] = 10'h191;
        mem[7] = 10'h201;
        mem[8] = 10'h0ba;
        mem[9] = 10'h159;
        mem[10] = 10'h36b;
        mem[11] = 10'h350;
        mem[12] = 10'h1fb;
        mem[13] = 10'h11f;
        mem[14] = 10'h33a;
        mem[15] = 10'h37f;
        mem[16] = 10'h1af;
        mem[17] = 10'h380;
        mem[18] = 10'h0ae;
        mem[19] = 10'h3c9;
        mem[20] = 10'h3c1;
        mem[21] = 10'h0dd;
        mem[22] = 10'h02d;
        mem[23] = 10'h16c;
        mem[24] = 10'h2d5;
        mem[25] = 10'h141;
        mem[26] = 10'h039;
        mem[27] = 10'h27e;
        mem[28] = 10'h315;
        mem[29] = 10'h109;
        mem[30] = 10'h234;
        mem[31] = 10'h241;
        mem[32] = 10'h335;
        mem[33] = 10'h39e;
        mem[34] = 10'h151;
        mem[35] = 10'h003;
        mem[36] = 10'h3d7;
        mem[37] = 10'h321;
        mem[38] = 10'h103;
        mem[39] = 10'h1bd;
        mem[40] = 10'h286;
        mem[41] = 10'h3df;
        mem[42] = 10'h1fd;
        mem[43] = 10'h2a0;
        mem[44] = 10'h35d;
        mem[45] = 10'h2ec;
        mem[46] = 10'h3a2;
        mem[47] = 10'h209;
        mem[48] = 10'h04a;
        mem[49] = 10'h079;
        mem[50] = 10'h165;
        mem[51] = 10'h01e;
        mem[52] = 10'h192;
        mem[53] = 10'h011;
        mem[54] = 10'h1d7;
        mem[55] = 10'h2e6;
        mem[56] = 10'h08b;
        mem[57] = 10'h161;
        mem[58] = 10'h397;
        mem[59] = 10'h19d;
        mem[60] = 10'h1ac;
        mem[61] = 10'h171;
        mem[62] = 10'h1e4;
        mem[63] = 10'h23d;
        mem[64] = 10'h046;
        mem[65] = 10'h3bf;
        mem[66] = 10'h1ed;
        mem[67] = 10'h12c;
        mem[68] = 10'h260;
        mem[69] = 10'h0ca;
        mem[70] = 10'h038;
        mem[71] = 10'h3b7;
        mem[72] = 10'h0ad;
        mem[73] = 10'h269;
        mem[74] = 10'h15f;
        mem[75] = 10'h085;
        mem[76] = 10'h263;
        mem[77] = 10'h123;
        mem[78] = 10'h3d1;
        mem[79] = 10'h162;
        mem[80] = 10'h1a9;
        mem[81] = 10'h1d8;
        mem[82] = 10'h3ce;
        mem[83] = 10'h2c2;
        mem[84] = 10'h096;
        mem[85] = 10'h235;
        mem[86] = 10'h32e;
        mem[87] = 10'h098;
        mem[88] = 10'h275;
        mem[89] = 10'h108;
        mem[90] = 10'h3c4;
        mem[91] = 10'h194;
        mem[92] = 10'h0bd;
        mem[93] = 10'h075;
        mem[94] = 10'h05b;
        mem[95] = 10'h0a1;
        mem[96] = 10'h13a;
        mem[97] = 10'h3f6;
        mem[98] = 10'h1cd;
        mem[99] = 10'h377;
        mem[100] = 10'h27b;
        mem[101] = 10'h35c;
        mem[102] = 10'h352;
        mem[103] = 10'h053;
        mem[104] = 10'h2fd;
        mem[105] = 10'h0a7;
        mem[106] = 10'h154;
        mem[107] = 10'h2a9;
        mem[108] = 10'h34a;
        mem[109] = 10'h238;
        mem[110] = 10'h1fc;
        mem[111] = 10'h1df;
        mem[112] = 10'h20f;
        mem[113] = 10'h3ac;
        mem[114] = 10'h03c;
        mem[115] = 10'h176;
        mem[116] = 10'h2c8;
        mem[117] = 10'h0ff;
        mem[118] = 10'h2ee;
        mem[119] = 10'h227;
        mem[120] = 10'h31f;
        mem[121] = 10'h3eb;
        mem[122] = 10'h131;
        mem[123] = 10'h290;
        mem[124] = 10'h1ef;
        mem[125] = 10'h38d;
        mem[126] = 10'h323;
        mem[127] = 10'h2eb;
        mem[128] = 10'h37a;
        mem[129] = 10'h18f;
        mem[130] = 10'h080;
        mem[131] = 10'h092;
        mem[132] = 10'h1da;
        mem[133] = 10'h1c3;
        mem[134] = 10'h12d;
        mem[135] = 10'h01d;
        mem[136] = 10'h239;
        mem[137] = 10'h3ba;
        mem[138] = 10'h399;
        mem[139] = 10'h2cc;
        mem[140] = 10'h115;
        mem[141] = 10'h2dd;
        mem[142] = 10'h040;
        mem[143] = 10'h088;
        mem[144] = 10'h170;
        mem[145] = 10'h26d;
        mem[146] = 10'h1f1;
        mem[147] = 10'h1a0;
        mem[148] = 10'h2b8;
        mem[149] = 10'h310;
        mem[150] = 10'h0b0;
        mem[151] = 10'h3d5;
        mem[152] = 10'h0c1;
        mem[153] = 10'h35f;
        mem[154] = 10'h0f3;
        mem[155] = 10'h3fb;
        mem[156] = 10'h0ee;
        mem[157] = 10'h158;
        mem[158] = 10'h300;
        mem[159] = 10'h03b;
        mem[160] = 10'h26a;
        mem[161] = 10'h3f2;
        mem[162] = 10'h272;
        mem[163] = 10'h3e7;
        mem[164] = 10'h2df;
        mem[165] = 10'h225;
        mem[166] = 10'h3b5;
        mem[167] = 10'h216;
        mem[168] = 10'h29a;
        mem[169] = 10'h1a7;
        mem[170] = 10'h230;
        mem[171] = 10'h1f7;
        mem[172] = 10'h247;
        mem[173] = 10'h0e8;
        mem[174] = 10'h200;
        mem[175] = 10'h089;
        mem[176] = 10'h1b1;
        mem[177] = 10'h364;
        mem[178] = 10'h250;
        mem[179] = 10'h1c5;
        mem[180] = 10'h135;
        mem[181] = 10'h13c;
        mem[182] = 10'h045;
        mem[183] = 10'h12e;
        mem[184] = 10'h3ab;
        mem[185] = 10'h274;
        mem[186] = 10'h39f;
        mem[187] = 10'h23c;
        mem[188] = 10'h18b;
        mem[189] = 10'h07a;
        mem[190] = 10'h386;
        mem[191] = 10'h266;
        mem[192] = 10'h1a3;
        mem[193] = 10'h06b;
        mem[194] = 10'h0bf;
        mem[195] = 10'h14f;
        mem[196] = 10'h308;
        mem[197] = 10'h35e;
        mem[198] = 10'h0d8;
        mem[199] = 10'h319;
        mem[200] = 10'h143;
        mem[201] = 10'h390;
        mem[202] = 10'h09e;
        mem[203] = 10'h385;
        mem[204] = 10'h21d;
        mem[205] = 10'h067;
        mem[206] = 10'h3f0;
        mem[207] = 10'h16d;
        mem[208] = 10'h355;
        mem[209] = 10'h3e5;
        mem[210] = 10'h2e4;
        mem[211] = 10'h177;
        mem[212] = 10'h3a4;
        mem[213] = 10'h24e;
        mem[214] = 10'h18a;
        mem[215] = 10'h31c;
        mem[216] = 10'h1f9;
        mem[217] = 10'h28a;
        mem[218] = 10'h3da;
        mem[219] = 10'h3d4;
        mem[220] = 10'h2bc;
        mem[221] = 10'h2ce;
        mem[222] = 10'h394;
        mem[223] = 10'h18c;
        mem[224] = 10'h343;
        mem[225] = 10'h20c;
        mem[226] = 10'h1a4;
        mem[227] = 10'h28c;
        mem[228] = 10'h1a1;
        mem[229] = 10'h05f;
        mem[230] = 10'h107;
        mem[231] = 10'h09a;
        mem[232] = 10'h39c;
        mem[233] = 10'h174;
        mem[234] = 10'h39b;
        mem[235] = 10'h3e3;
        mem[236] = 10'h04b;
        mem[237] = 10'h1e6;
        mem[238] = 10'h010;
        mem[239] = 10'h21e;
        mem[240] = 10'h059;
        mem[241] = 10'h0de;
        mem[242] = 10'h39a;
        mem[243] = 10'h3fc;
        mem[244] = 10'h2f4;
        mem[245] = 10'h000;
        mem[246] = 10'h1ba;
        mem[247] = 10'h24d;
        mem[248] = 10'h268;
        mem[249] = 10'h28e;
        mem[250] = 10'h2b6;
        mem[251] = 10'h17c;
        mem[252] = 10'h102;
        mem[253] = 10'h071;
        mem[254] = 10'h055;
        mem[255] = 10'h023;
        mem[256] = 10'h220;
        mem[257] = 10'h281;
        mem[258] = 10'h1ae;
        mem[259] = 10'h1fa;
        mem[260] = 10'h1dc;
        mem[261] = 10'h1c1;
        mem[262] = 10'h0ea;
        mem[263] = 10'h1dd;
        mem[264] = 10'h33e;
        mem[265] = 10'h25a;
        mem[266] = 10'h0ce;
        mem[267] = 10'h093;
        mem[268] = 10'h140;
        mem[269] = 10'h150;
        mem[270] = 10'h188;
        mem[271] = 10'h169;
        mem[272] = 10'h344;
        mem[273] = 10'h0b8;
        mem[274] = 10'h189;
        mem[275] = 10'h0d9;
        mem[276] = 10'h16b;
        mem[277] = 10'h070;
        mem[278] = 10'h2fc;
        mem[279] = 10'h1a2;
        mem[280] = 10'h1b4;
        mem[281] = 10'h178;
        mem[282] = 10'h2d7;
        mem[283] = 10'h047;
        mem[284] = 10'h1c6;
        mem[285] = 10'h2c9;
        mem[286] = 10'h01a;
        mem[287] = 10'h257;
        mem[288] = 10'h2e1;
        mem[289] = 10'h16e;
        mem[290] = 10'h0bb;
        mem[291] = 10'h255;
        mem[292] = 10'h23b;
        mem[293] = 10'h183;
        mem[294] = 10'h3db;
        mem[295] = 10'h07f;
        mem[296] = 10'h16a;
        mem[297] = 10'h298;
        mem[298] = 10'h15b;
        mem[299] = 10'h0e3;
        mem[300] = 10'h312;
        mem[301] = 10'h2d6;
        mem[302] = 10'h2d3;
        mem[303] = 10'h2a7;
        mem[304] = 10'h001;
        mem[305] = 10'h212;
        mem[306] = 10'h1db;
        mem[307] = 10'h0e4;
        mem[308] = 10'h016;
        mem[309] = 10'h042;
        mem[310] = 10'h2f9;
        mem[311] = 10'h357;
        mem[312] = 10'h0fe;
        mem[313] = 10'h3ad;
        mem[314] = 10'h396;
        mem[315] = 10'h05a;
        mem[316] = 10'h3de;
        mem[317] = 10'h187;
        mem[318] = 10'h083;
        mem[319] = 10'h2f3;
        mem[320] = 10'h336;
        mem[321] = 10'h2f5;
        mem[322] = 10'h1e5;
        mem[323] = 10'h237;
        mem[324] = 10'h0d0;
        mem[325] = 10'h122;
        mem[326] = 10'h02c;
        mem[327] = 10'h2e7;
        mem[328] = 10'h18e;
        mem[329] = 10'h06f;
        mem[330] = 10'h1e8;
        mem[331] = 10'h13e;
        mem[332] = 10'h236;
        mem[333] = 10'h1b6;
        mem[334] = 10'h3a8;
        mem[335] = 10'h366;
        mem[336] = 10'h2d2;
        mem[337] = 10'h2cb;
        mem[338] = 10'h0c8;
        mem[339] = 10'h1b2;
        mem[340] = 10'h19e;
        mem[341] = 10'h121;
        mem[342] = 10'h2e0;
        mem[343] = 10'h2c7;
        mem[344] = 10'h284;
        mem[345] = 10'h1d2;
        mem[346] = 10'h2ad;
        mem[347] = 10'h113;
        mem[348] = 10'h27d;
        mem[349] = 10'h2ed;
        mem[350] = 10'h1aa;
        mem[351] = 10'h0f0;
        mem[352] = 10'h025;
        mem[353] = 10'h3b9;
        mem[354] = 10'h379;
        mem[355] = 10'h07e;
        mem[356] = 10'h2c1;
        mem[357] = 10'h14e;
        mem[358] = 10'h3cd;
        mem[359] = 10'h112;
        mem[360] = 10'h0a9;
        mem[361] = 10'h3f5;
        mem[362] = 10'h243;
        mem[363] = 10'h196;
        mem[364] = 10'h2e9;
        mem[365] = 10'h04f;
        mem[366] = 10'h1c4;
        mem[367] = 10'h26f;
        mem[368] = 10'h3f3;
        mem[369] = 10'h0f2;
        mem[370] = 10'h127;
        mem[371] = 10'h17a;
        mem[372] = 10'h0d6;
        mem[373] = 10'h0d2;
        mem[374] = 10'h3a1;
        mem[375] = 10'h0cb;
        mem[376] = 10'h3c7;
        mem[377] = 10'h1b3;
        mem[378] = 10'h181;
        mem[379] = 10'h1f4;
        mem[380] = 10'h197;
        mem[381] = 10'h0c7;
        mem[382] = 10'h12b;
        mem[383] = 10'h0d1;
        mem[384] = 10'h152;
        mem[385] = 10'h288;
        mem[386] = 10'h14a;
        mem[387] = 10'h3f7;
        mem[388] = 10'h251;
        mem[389] = 10'h26b;
        mem[390] = 10'h228;
        mem[391] = 10'h322;
        mem[392] = 10'h3af;
        mem[393] = 10'h03f;
        mem[394] = 10'h3be;
        mem[395] = 10'h044;
        mem[396] = 10'h2cd;
        mem[397] = 10'h3e2;
        mem[398] = 10'h3bd;
        mem[399] = 10'h1bf;
        mem[400] = 10'h15c;
        mem[401] = 10'h273;
        mem[402] = 10'h0af;
        mem[403] = 10'h287;
        mem[404] = 10'h305;
        mem[405] = 10'h3ae;
        mem[406] = 10'h324;
        mem[407] = 10'h175;
        mem[408] = 10'h0f9;
        mem[409] = 10'h29e;
        mem[410] = 10'h28b;
        mem[411] = 10'h1e9;
        mem[412] = 10'h34c;
        mem[413] = 10'h128;
        mem[414] = 10'h11e;
        mem[415] = 10'h09f;
        mem[416] = 10'h27f;
        mem[417] = 10'h198;
        mem[418] = 10'h0b7;
        mem[419] = 10'h1d0;
        mem[420] = 10'h278;
        mem[421] = 10'h020;
        mem[422] = 10'h39d;
        mem[423] = 10'h2be;
        mem[424] = 10'h069;
        mem[425] = 10'h2ba;
        mem[426] = 10'h087;
        mem[427] = 10'h168;
        mem[428] = 10'h334;
        mem[429] = 10'h017;
        mem[430] = 10'h095;
        mem[431] = 10'h2c6;
        mem[432] = 10'h01b;
        mem[433] = 10'h13d;
        mem[434] = 10'h20b;
        mem[435] = 10'h370;
        mem[436] = 10'h1c9;
        mem[437] = 10'h3c3;
        mem[438] = 10'h37c;
        mem[439] = 10'h048;
        mem[440] = 10'h0db;
        mem[441] = 10'h1a8;
        mem[442] = 10'h2b7;
        mem[443] = 10'h362;
        mem[444] = 10'h389;
        mem[445] = 10'h28f;
        mem[446] = 10'h17f;
        mem[447] = 10'h0c4;
        mem[448] = 10'h34d;
        mem[449] = 10'h211;
        mem[450] = 10'h0a2;
        mem[451] = 10'h10c;
        mem[452] = 10'h244;
        mem[453] = 10'h307;
        mem[454] = 10'h374;
        mem[455] = 10'h05d;
        mem[456] = 10'h339;
        mem[457] = 10'h2b0;
        mem[458] = 10'h378;
        mem[459] = 10'h073;
        mem[460] = 10'h144;
        mem[461] = 10'h056;
        mem[462] = 10'h118;
        mem[463] = 10'h10e;
        mem[464] = 10'h057;
        mem[465] = 10'h19c;
        mem[466] = 10'h34f;
        mem[467] = 10'h28d;
        mem[468] = 10'h17b;
        mem[469] = 10'h361;
        mem[470] = 10'h180;
        mem[471] = 10'h10b;
        mem[472] = 10'h106;
        mem[473] = 10'h293;
        mem[474] = 10'h02b;
        mem[475] = 10'h294;
        mem[476] = 10'h0c5;
        mem[477] = 10'h2a8;
        mem[478] = 10'h218;
        mem[479] = 10'h110;
        mem[480] = 10'h10f;
        mem[481] = 10'h08f;
        mem[482] = 10'h149;
        mem[483] = 10'h398;
        mem[484] = 10'h330;
        mem[485] = 10'h20d;
        mem[486] = 10'h30e;
        mem[487] = 10'h265;
        mem[488] = 10'h254;
        mem[489] = 10'h33b;
        mem[490] = 10'h25f;
        mem[491] = 10'h291;
        mem[492] = 10'h0e5;
        mem[493] = 10'h327;
        mem[494] = 10'h022;
        mem[495] = 10'h14c;
        mem[496] = 10'h014;
        mem[497] = 10'h17e;
        mem[498] = 10'h086;
        mem[499] = 10'h1b5;
        mem[500] = 10'h1c0;
        mem[501] = 10'h0cc;
        mem[502] = 10'h3f8;
        mem[503] = 10'h204;
        mem[504] = 10'h0b9;
        mem[505] = 10'h354;
        mem[506] = 10'h31d;
        mem[507] = 10'h060;
        mem[508] = 10'h147;
        mem[509] = 10'h3ef;
        mem[510] = 10'h054;
        mem[511] = 10'h232;
        mem[512] = 10'h19b;
        mem[513] = 10'h0d4;
        mem[514] = 10'h076;
        mem[515] = 10'h07b;
        mem[516] = 10'h2d9;
        mem[517] = 10'h1e1;
        mem[518] = 10'h31b;
        mem[519] = 10'h316;
        mem[520] = 10'h2af;
        mem[521] = 10'h215;
        mem[522] = 10'h1f8;
        mem[523] = 10'h217;
        mem[524] = 10'h136;
        mem[525] = 10'h2d8;
        mem[526] = 10'h116;
        mem[527] = 10'h08d;
        mem[528] = 10'h2b1;
        mem[529] = 10'h21c;
        mem[530] = 10'h12f;
        mem[531] = 10'h077;
        mem[532] = 10'h262;
        mem[533] = 10'h372;
        mem[534] = 10'h138;
        mem[535] = 10'h369;
        mem[536] = 10'h393;
        mem[537] = 10'h10d;
        mem[538] = 10'h0ab;
        mem[539] = 10'h1d6;
        mem[540] = 10'h1eb;
        mem[541] = 10'h09b;
        mem[542] = 10'h156;
        mem[543] = 10'h1a6;
        mem[544] = 10'h37e;
        mem[545] = 10'h302;
        mem[546] = 10'h1f0;
        mem[547] = 10'h249;
        mem[548] = 10'h3d8;
        mem[549] = 10'h0cd;
        mem[550] = 10'h2e5;
        mem[551] = 10'h0f4;
        mem[552] = 10'h356;
        mem[553] = 10'h30f;
        mem[554] = 10'h0c3;
        mem[555] = 10'h25d;
        mem[556] = 10'h30d;
        mem[557] = 10'h006;
        mem[558] = 10'h13f;
        mem[559] = 10'h384;
        mem[560] = 10'h311;
        mem[561] = 10'h050;
        mem[562] = 10'h2cf;
        mem[563] = 10'h3ca;
        mem[564] = 10'h27a;
        mem[565] = 10'h373;
        mem[566] = 10'h030;
        mem[567] = 10'h29c;
        mem[568] = 10'h114;
        mem[569] = 10'h2ae;
        mem[570] = 10'h2a1;
        mem[571] = 10'h277;
        mem[572] = 10'h018;
        mem[573] = 10'h1ee;
        mem[574] = 10'h231;
        mem[575] = 10'h3cc;
        mem[576] = 10'h0a8;
        mem[577] = 10'h3e0;
        mem[578] = 10'h2b4;
        mem[579] = 10'h341;
        mem[580] = 10'h021;
        mem[581] = 10'h0a0;
        mem[582] = 10'h2c0;
        mem[583] = 10'h34b;
        mem[584] = 10'h376;
        mem[585] = 10'h0c0;
        mem[586] = 10'h329;
        mem[587] = 10'h347;
        mem[588] = 10'h1ca;
        mem[589] = 10'h3fe;
        mem[590] = 10'h224;
        mem[591] = 10'h233;
        mem[592] = 10'h304;
        mem[593] = 10'h383;
        mem[594] = 10'h29f;
        mem[595] = 10'h19a;
        mem[596] = 10'h1f5;
        mem[597] = 10'h0e6;
        mem[598] = 10'h11a;
        mem[599] = 10'h345;
        mem[600] = 10'h205;
        mem[601] = 10'h005;
        mem[602] = 10'h3aa;
        mem[603] = 10'h3f4;
        mem[604] = 10'h229;
        mem[605] = 10'h2d0;
        mem[606] = 10'h0fb;
        mem[607] = 10'h296;
        mem[608] = 10'h024;
        mem[609] = 10'h2b3;
        mem[610] = 10'h03a;
        mem[611] = 10'h338;
        mem[612] = 10'h3a5;
        mem[613] = 10'h11d;
        mem[614] = 10'h270;
        mem[615] = 10'h2ef;
        mem[616] = 10'h317;
        mem[617] = 10'h0aa;
        mem[618] = 10'h019;
        mem[619] = 10'h2bb;
        mem[620] = 10'h1d5;
        mem[621] = 10'h1ec;
        mem[622] = 10'h04e;
        mem[623] = 10'h353;
        mem[624] = 10'h049;
        mem[625] = 10'h22e;
        mem[626] = 10'h371;
        mem[627] = 10'h125;
        mem[628] = 10'h3ee;
        mem[629] = 10'h30b;
        mem[630] = 10'h2a5;
        mem[631] = 10'h282;
        mem[632] = 10'h193;
        mem[633] = 10'h2e3;
        mem[634] = 10'h035;
        mem[635] = 10'h3d6;
        mem[636] = 10'h142;
        mem[637] = 10'h3a0;
        mem[638] = 10'h1ff;
        mem[639] = 10'h26e;
        mem[640] = 10'h32d;
        mem[641] = 10'h395;
        mem[642] = 10'h360;
        mem[643] = 10'h23a;
        mem[644] = 10'h063;
        mem[645] = 10'h35a;
        mem[646] = 10'h223;
        mem[647] = 10'h3ed;
        mem[648] = 10'h1ea;
        mem[649] = 10'h289;
        mem[650] = 10'h0be;
        mem[651] = 10'h099;
        mem[652] = 10'h1ad;
        mem[653] = 10'h276;
        mem[654] = 10'h3e8;
        mem[655] = 10'h245;
        mem[656] = 10'h0c6;
        mem[657] = 10'h325;
        mem[658] = 10'h253;
        mem[659] = 10'h210;
        mem[660] = 10'h0ac;
        mem[661] = 10'h332;
        mem[662] = 10'h3d9;
        mem[663] = 10'h23e;
        mem[664] = 10'h213;
        mem[665] = 10'h1d9;
        mem[666] = 10'h148;
        mem[667] = 10'h3c8;
        mem[668] = 10'h034;
        mem[669] = 10'h24a;
        mem[670] = 10'h31a;
        mem[671] = 10'h1e7;
        mem[672] = 10'h004;
        mem[673] = 10'h2d4;
        mem[674] = 10'h0ef;
        mem[675] = 10'h061;
        mem[676] = 10'h21a;
        mem[677] = 10'h101;
        mem[678] = 10'h1e3;
        mem[679] = 10'h358;
        mem[680] = 10'h0a6;
        mem[681] = 10'h081;
        mem[682] = 10'h29b;
        mem[683] = 10'h359;
        mem[684] = 10'h303;
        mem[685] = 10'h27c;
        mem[686] = 10'h221;
        mem[687] = 10'h22b;
        mem[688] = 10'h2e8;
        mem[689] = 10'h2da;
        mem[690] = 10'h32a;
        mem[691] = 10'h1b9;
        mem[692] = 10'h16f;
        mem[693] = 10'h133;
        mem[694] = 10'h02e;
        mem[695] = 10'h381;
        mem[696] = 10'h026;
        mem[697] = 10'h1f2;
        mem[698] = 10'h134;
        mem[699] = 10'h283;
        mem[700] = 10'h14d;
        mem[701] = 10'h219;
        mem[702] = 10'h3a7;
        mem[703] = 10'h29d;
        mem[704] = 10'h01f;
        mem[705] = 10'h1bc;
        mem[706] = 10'h06c;
        mem[707] = 10'h22d;
        mem[708] = 10'h068;
        mem[709] = 10'h38a;
        mem[710] = 10'h1de;
        mem[711] = 10'h21f;
        mem[712] = 10'h2a3;
        mem[713] = 10'h0e9;
        mem[714] = 10'h12a;
        mem[715] = 10'h09c;
        mem[716] = 10'h097;
        mem[717] = 10'h1c2;
        mem[718] = 10'h0b3;
        mem[719] = 10'h06a;
        mem[720] = 10'h35b;
        mem[721] = 10'h111;
        mem[722] = 10'h202;
        mem[723] = 10'h348;
        mem[724] = 10'h15a;
        mem[725] = 10'h094;
        mem[726] = 10'h1cf;
        mem[727] = 10'h267;
        mem[728] = 10'h153;
        mem[729] = 10'h08c;
        mem[730] = 10'h203;
        mem[731] = 10'h041;
        mem[732] = 10'h160;
        mem[733] = 10'h349;
        mem[734] = 10'h032;
        mem[735] = 10'h2c5;
        mem[736] = 10'h3c5;
        mem[737] = 10'h3dd;
        mem[738] = 10'h084;
        mem[739] = 10'h06d;
        mem[740] = 10'h2ea;
        mem[741] = 10'h3f1;
        mem[742] = 10'h0dc;
        mem[743] = 10'h34e;
        mem[744] = 10'h363;
        mem[745] = 10'h02a;
        mem[746] = 10'h365;
        mem[747] = 10'h1e0;
        mem[748] = 10'h0e2;
        mem[749] = 10'h3ff;
        mem[750] = 10'h246;
        mem[751] = 10'h090;
        mem[752] = 10'h13b;
        mem[753] = 10'h3d0;
        mem[754] = 10'h0ec;
        mem[755] = 10'h013;
        mem[756] = 10'h027;
        mem[757] = 10'h392;
        mem[758] = 10'h04c;
        mem[759] = 10'h07d;
        mem[760] = 10'h066;
        mem[761] = 10'h388;
        mem[762] = 10'h3e4;
        mem[763] = 10'h1c7;
        mem[764] = 10'h32b;
        mem[765] = 10'h0a4;
        mem[766] = 10'h15d;
        mem[767] = 10'h002;
        mem[768] = 10'h2ca;
        mem[769] = 10'h2f2;
        mem[770] = 10'h172;
        mem[771] = 10'h078;
        mem[772] = 10'h182;
        mem[773] = 10'h37b;
        mem[774] = 10'h2f0;
        mem[775] = 10'h1b0;
        mem[776] = 10'h0d5;
        mem[777] = 10'h0d3;
        mem[778] = 10'h375;
        mem[779] = 10'h346;
        mem[780] = 10'h38e;
        mem[781] = 10'h3b8;
        mem[782] = 10'h280;
        mem[783] = 10'h02f;
        mem[784] = 10'h1a5;
        mem[785] = 10'h32f;
        mem[786] = 10'h173;
        mem[787] = 10'h185;
        mem[788] = 10'h2f1;
        mem[789] = 10'h164;
        mem[790] = 10'h2e2;
        mem[791] = 10'h1bb;
        mem[792] = 10'h285;
        mem[793] = 10'h297;
        mem[794] = 10'h342;
        mem[795] = 10'h05c;
        mem[796] = 10'h146;
        mem[797] = 10'h1ce;
        mem[798] = 10'h0c2;
        mem[799] = 10'h36d;
        mem[800] = 10'h074;
        mem[801] = 10'h3fa;
        mem[802] = 10'h258;
        mem[803] = 10'h0e0;
        mem[804] = 10'h11c;
        mem[805] = 10'h166;
        mem[806] = 10'h2ff;
        mem[807] = 10'h37d;
        mem[808] = 10'h208;
        mem[809] = 10'h0e1;
        mem[810] = 10'h1ab;
        mem[811] = 10'h17d;
        mem[812] = 10'h00a;
        mem[813] = 10'h252;
        mem[814] = 10'h33c;
        mem[815] = 10'h3ea;
        mem[816] = 10'h139;
        mem[817] = 10'h261;
        mem[818] = 10'h3b0;
        mem[819] = 10'h31e;
        mem[820] = 10'h214;
        mem[821] = 10'h0df;
        mem[822] = 10'h3b6;
        mem[823] = 10'h2db;
        mem[824] = 10'h22f;
        mem[825] = 10'h2b9;
        mem[826] = 10'h2dc;
        mem[827] = 10'h179;
        mem[828] = 10'h008;
        mem[829] = 10'h2f6;
        mem[830] = 10'h1b7;
        mem[831] = 10'h117;
        mem[832] = 10'h3dc;
        mem[833] = 10'h33f;
        mem[834] = 10'h0b6;
        mem[835] = 10'h105;
        mem[836] = 10'h11b;
        mem[837] = 10'h0bc;
        mem[838] = 10'h01c;
        mem[839] = 10'h2d1;
        mem[840] = 10'h00d;
        mem[841] = 10'h248;
        mem[842] = 10'h22a;
        mem[843] = 10'h0fa;
        mem[844] = 10'h0e7;
        mem[845] = 10'h36e;
        mem[846] = 10'h00b;
        mem[847] = 10'h2aa;
        mem[848] = 10'h0f6;
        mem[849] = 10'h2fa;
        mem[850] = 10'h2f7;
        mem[851] = 10'h0b4;
        mem[852] = 10'h2b2;
        mem[853] = 10'h119;
        mem[854] = 10'h037;
        mem[855] = 10'h043;
        mem[856] = 10'h1b8;
        mem[857] = 10'h036;
        mem[858] = 10'h3b4;
        mem[859] = 10'h26c;
        mem[860] = 10'h3e1;
        mem[861] = 10'h259;
        mem[862] = 10'h0ed;
        mem[863] = 10'h3b3;
        mem[864] = 10'h3d3;
        mem[865] = 10'h3c6;
        mem[866] = 10'h130;
        mem[867] = 10'h06e;
        mem[868] = 10'h318;
        mem[869] = 10'h0a3;
        mem[870] = 10'h3b2;
        mem[871] = 10'h23f;
        mem[872] = 10'h167;
        mem[873] = 10'h120;
        mem[874] = 10'h129;
        mem[875] = 10'h306;
        mem[876] = 10'h100;
        mem[877] = 10'h299;
        mem[878] = 10'h1cc;
        mem[879] = 10'h2bd;
        mem[880] = 10'h0f7;
        mem[881] = 10'h226;
        mem[882] = 10'h155;
        mem[883] = 10'h3bc;
        mem[884] = 10'h314;
        mem[885] = 10'h3c2;
        mem[886] = 10'h25c;
        mem[887] = 10'h3a9;
        mem[888] = 10'h0d7;
        mem[889] = 10'h07c;
        mem[890] = 10'h382;
        mem[891] = 10'h3cf;
        mem[892] = 10'h295;
        mem[893] = 10'h3a3;
        mem[894] = 10'h072;
        mem[895] = 10'h029;
        mem[896] = 10'h32c;
        mem[897] = 10'h391;
        mem[898] = 10'h1d4;
        mem[899] = 10'h00f;
        mem[900] = 10'h1f6;
        mem[901] = 10'h2a6;
        mem[902] = 10'h1c8;
        mem[903] = 10'h3f9;
        mem[904] = 10'h0b5;
        mem[905] = 10'h340;
        mem[906] = 10'h292;
        mem[907] = 10'h012;
        mem[908] = 10'h2b5;
        mem[909] = 10'h206;
        mem[910] = 10'h328;
        mem[911] = 10'h21b;
        mem[912] = 10'h22c;
        mem[913] = 10'h2ab;
        mem[914] = 10'h082;
        mem[915] = 10'h326;
        mem[916] = 10'h0f1;
        mem[917] = 10'h3d2;
        mem[918] = 10'h3e6;
        mem[919] = 10'h132;
        mem[920] = 10'h0da;
        mem[921] = 10'h256;
        mem[922] = 10'h14b;
        mem[923] = 10'h051;
        mem[924] = 10'h00c;
        mem[925] = 10'h2fb;
        mem[926] = 10'h20a;
        mem[927] = 10'h368;
        mem[928] = 10'h38f;
        mem[929] = 10'h03e;
        mem[930] = 10'h25e;
        mem[931] = 10'h190;
        mem[932] = 10'h091;
        mem[933] = 10'h18d;
        mem[934] = 10'h24b;
        mem[935] = 10'h367;
        mem[936] = 10'h38c;
        mem[937] = 10'h3c0;
        mem[938] = 10'h052;
        mem[939] = 10'h313;
        mem[940] = 10'h279;
        mem[941] = 10'h09d;
        mem[942] = 10'h2f8;
        mem[943] = 10'h163;
        mem[944] = 10'h301;
        mem[945] = 10'h1d3;
        mem[946] = 10'h242;
        mem[947] = 10'h3cb;
        mem[948] = 10'h240;
        mem[949] = 10'h186;
        mem[950] = 10'h320;
        mem[951] = 10'h25b;
        mem[952] = 10'h0b1;
        mem[953] = 10'h145;
        mem[954] = 10'h0a5;
        mem[955] = 10'h331;
        mem[956] = 10'h19f;
        mem[957] = 10'h1d1;
        mem[958] = 10'h10a;
        mem[959] = 10'h309;
        mem[960] = 10'h2a4;
        mem[961] = 10'h064;
        mem[962] = 10'h36c;
        mem[963] = 10'h04d;
        mem[964] = 10'h03d;
        mem[965] = 10'h0b2;
        mem[966] = 10'h2c3;
        mem[967] = 10'h031;
        mem[968] = 10'h337;
        mem[969] = 10'h3a6;
        mem[970] = 10'h0c9;
        mem[971] = 10'h264;
        mem[972] = 10'h062;
        mem[973] = 10'h387;
        mem[974] = 10'h24f;
        mem[975] = 10'h3ec;
        mem[976] = 10'h2ac;
        mem[977] = 10'h1be;
        mem[978] = 10'h1cb;
        mem[979] = 10'h184;
        mem[980] = 10'h271;
        mem[981] = 10'h028;
        mem[982] = 10'h1e2;
        mem[983] = 10'h222;
        mem[984] = 10'h1f3;
        mem[985] = 10'h36a;
        mem[986] = 10'h333;
        mem[987] = 10'h058;
        mem[988] = 10'h1fe;
        mem[989] = 10'h2bf;
        mem[990] = 10'h2de;
        mem[991] = 10'h30a;
        mem[992] = 10'h24c;
        mem[993] = 10'h2c4;
        mem[994] = 10'h33d;
        mem[995] = 10'h065;
        mem[996] = 10'h20e;
        mem[997] = 10'h033;
        mem[998] = 10'h007;
        mem[999] = 10'h157;
        mem[1000] = 10'h124;
        mem[1001] = 10'h199;
        mem[1002] = 10'h2a2;
        mem[1003] = 10'h3b1;
        mem[1004] = 10'h351;
        mem[1005] = 10'h0fd;
        mem[1006] = 10'h00e;
        mem[1007] = 10'h08e;
        mem[1008] = 10'h0f5;
        mem[1009] = 10'h05e;
        mem[1010] = 10'h015;
        mem[1011] = 10'h15e;
        mem[1012] = 10'h0fc;
        mem[1013] = 10'h0cf;
        mem[1014] = 10'h3bb;
        mem[1015] = 10'h137;
        mem[1016] = 10'h08a;
        mem[1017] = 10'h3e9;
        mem[1018] = 10'h30c;
        mem[1019] = 10'h195;
        mem[1020] = 10'h0eb;
        mem[1021] = 10'h104;
        mem[1022] = 10'h126;
        mem[1023] = 10'h009;
    end
endmodule

module odo_sbox_large9(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h3a3;
        mem[1] = 10'h2b1;
        mem[2] = 10'h243;
        mem[3] = 10'h1b5;
        mem[4] = 10'h12c;
        mem[5] = 10'h004;
        mem[6] = 10'h3c0;
        mem[7] = 10'h3a6;
        mem[8] = 10'h2cd;
        mem[9] = 10'h364;
        mem[10] = 10'h0e0;
        mem[11] = 10'h3cf;
        mem[12] = 10'h21a;
        mem[13] = 10'h15f;
        mem[14] = 10'h0a0;
        mem[15] = 10'h204;
        mem[16] = 10'h062;
        mem[17] = 10'h135;
        mem[18] = 10'h356;
        mem[19] = 10'h274;
        mem[20] = 10'h2be;
        mem[21] = 10'h337;
        mem[22] = 10'h177;
        mem[23] = 10'h016;
        mem[24] = 10'h1b0;
        mem[25] = 10'h354;
        mem[26] = 10'h339;
        mem[27] = 10'h256;
        mem[28] = 10'h2c5;
        mem[29] = 10'h30c;
        mem[30] = 10'h312;
        mem[31] = 10'h154;
        mem[32] = 10'h3c7;
        mem[33] = 10'h06b;
        mem[34] = 10'h09b;
        mem[35] = 10'h388;
        mem[36] = 10'h1a3;
        mem[37] = 10'h014;
        mem[38] = 10'h0f4;
        mem[39] = 10'h241;
        mem[40] = 10'h2c4;
        mem[41] = 10'h171;
        mem[42] = 10'h1ce;
        mem[43] = 10'h303;
        mem[44] = 10'h335;
        mem[45] = 10'h1b1;
        mem[46] = 10'h2db;
        mem[47] = 10'h333;
        mem[48] = 10'h317;
        mem[49] = 10'h083;
        mem[50] = 10'h039;
        mem[51] = 10'h389;
        mem[52] = 10'h036;
        mem[53] = 10'h08a;
        mem[54] = 10'h078;
        mem[55] = 10'h071;
        mem[56] = 10'h1c3;
        mem[57] = 10'h060;
        mem[58] = 10'h14f;
        mem[59] = 10'h28e;
        mem[60] = 10'h168;
        mem[61] = 10'h010;
        mem[62] = 10'h151;
        mem[63] = 10'h259;
        mem[64] = 10'h017;
        mem[65] = 10'h382;
        mem[66] = 10'h2d8;
        mem[67] = 10'h10e;
        mem[68] = 10'h340;
        mem[69] = 10'h0e1;
        mem[70] = 10'h08c;
        mem[71] = 10'h104;
        mem[72] = 10'h279;
        mem[73] = 10'h305;
        mem[74] = 10'h2ba;
        mem[75] = 10'h0de;
        mem[76] = 10'h1f9;
        mem[77] = 10'h36a;
        mem[78] = 10'h103;
        mem[79] = 10'h0a8;
        mem[80] = 10'h267;
        mem[81] = 10'h0b8;
        mem[82] = 10'h12a;
        mem[83] = 10'h184;
        mem[84] = 10'h2da;
        mem[85] = 10'h3bf;
        mem[86] = 10'h0fb;
        mem[87] = 10'h254;
        mem[88] = 10'h113;
        mem[89] = 10'h234;
        mem[90] = 10'h36b;
        mem[91] = 10'h2f5;
        mem[92] = 10'h304;
        mem[93] = 10'h2ee;
        mem[94] = 10'h150;
        mem[95] = 10'h061;
        mem[96] = 10'h023;
        mem[97] = 10'h159;
        mem[98] = 10'h23f;
        mem[99] = 10'h237;
        mem[100] = 10'h05a;
        mem[101] = 10'h027;
        mem[102] = 10'h346;
        mem[103] = 10'h349;
        mem[104] = 10'h381;
        mem[105] = 10'h141;
        mem[106] = 10'h2e6;
        mem[107] = 10'h191;
        mem[108] = 10'h1a7;
        mem[109] = 10'h0ec;
        mem[110] = 10'h280;
        mem[111] = 10'h2bd;
        mem[112] = 10'h3b9;
        mem[113] = 10'h3cd;
        mem[114] = 10'h212;
        mem[115] = 10'h3ca;
        mem[116] = 10'h3e7;
        mem[117] = 10'h288;
        mem[118] = 10'h0af;
        mem[119] = 10'h39e;
        mem[120] = 10'h248;
        mem[121] = 10'h253;
        mem[122] = 10'h041;
        mem[123] = 10'h160;
        mem[124] = 10'h109;
        mem[125] = 10'h363;
        mem[126] = 10'h29b;
        mem[127] = 10'h278;
        mem[128] = 10'h327;
        mem[129] = 10'h158;
        mem[130] = 10'h37b;
        mem[131] = 10'h32a;
        mem[132] = 10'h322;
        mem[133] = 10'h1d8;
        mem[134] = 10'h34f;
        mem[135] = 10'h2c2;
        mem[136] = 10'h2d2;
        mem[137] = 10'h1e3;
        mem[138] = 10'h2ec;
        mem[139] = 10'h07c;
        mem[140] = 10'h043;
        mem[141] = 10'h0ea;
        mem[142] = 10'h198;
        mem[143] = 10'h180;
        mem[144] = 10'h37e;
        mem[145] = 10'h28d;
        mem[146] = 10'h034;
        mem[147] = 10'h0dd;
        mem[148] = 10'h0ab;
        mem[149] = 10'h33d;
        mem[150] = 10'h0a3;
        mem[151] = 10'h0ac;
        mem[152] = 10'h3b4;
        mem[153] = 10'h2b8;
        mem[154] = 10'h01b;
        mem[155] = 10'h11a;
        mem[156] = 10'h219;
        mem[157] = 10'h045;
        mem[158] = 10'h10a;
        mem[159] = 10'h139;
        mem[160] = 10'h136;
        mem[161] = 10'h2bc;
        mem[162] = 10'h0e2;
        mem[163] = 10'h36d;
        mem[164] = 10'h0f1;
        mem[165] = 10'h03c;
        mem[166] = 10'h3c1;
        mem[167] = 10'h226;
        mem[168] = 10'h0c8;
        mem[169] = 10'h162;
        mem[170] = 10'h32c;
        mem[171] = 10'h3b2;
        mem[172] = 10'h125;
        mem[173] = 10'h1a9;
        mem[174] = 10'h112;
        mem[175] = 10'h371;
        mem[176] = 10'h27a;
        mem[177] = 10'h03a;
        mem[178] = 10'h245;
        mem[179] = 10'h133;
        mem[180] = 10'h39a;
        mem[181] = 10'h011;
        mem[182] = 10'h222;
        mem[183] = 10'h2b3;
        mem[184] = 10'h0f8;
        mem[185] = 10'h244;
        mem[186] = 10'h3bb;
        mem[187] = 10'h28c;
        mem[188] = 10'h147;
        mem[189] = 10'h343;
        mem[190] = 10'h2a4;
        mem[191] = 10'h31e;
        mem[192] = 10'h143;
        mem[193] = 10'h301;
        mem[194] = 10'h2d0;
        mem[195] = 10'h3d6;
        mem[196] = 10'h086;
        mem[197] = 10'h203;
        mem[198] = 10'h208;
        mem[199] = 10'h1ae;
        mem[200] = 10'h39f;
        mem[201] = 10'h063;
        mem[202] = 10'h106;
        mem[203] = 10'h36c;
        mem[204] = 10'h2e9;
        mem[205] = 10'h19d;
        mem[206] = 10'h277;
        mem[207] = 10'h048;
        mem[208] = 10'h14c;
        mem[209] = 10'h1f5;
        mem[210] = 10'h372;
        mem[211] = 10'h3ed;
        mem[212] = 10'h270;
        mem[213] = 10'h19c;
        mem[214] = 10'h38d;
        mem[215] = 10'h05c;
        mem[216] = 10'h264;
        mem[217] = 10'h157;
        mem[218] = 10'h134;
        mem[219] = 10'h2a2;
        mem[220] = 10'h117;
        mem[221] = 10'h3d1;
        mem[222] = 10'h3fe;
        mem[223] = 10'h3f7;
        mem[224] = 10'h194;
        mem[225] = 10'h2e2;
        mem[226] = 10'h2f8;
        mem[227] = 10'h2d5;
        mem[228] = 10'h1c7;
        mem[229] = 10'h17e;
        mem[230] = 10'h137;
        mem[231] = 10'h0ba;
        mem[232] = 10'h37d;
        mem[233] = 10'h26a;
        mem[234] = 10'h1ff;
        mem[235] = 10'h02c;
        mem[236] = 10'h1bd;
        mem[237] = 10'h2de;
        mem[238] = 10'h20b;
        mem[239] = 10'h20e;
        mem[240] = 10'h351;
        mem[241] = 10'h18e;
        mem[242] = 10'h26c;
        mem[243] = 10'h1c9;
        mem[244] = 10'h090;
        mem[245] = 10'h072;
        mem[246] = 10'h1a4;
        mem[247] = 10'h146;
        mem[248] = 10'h0d7;
        mem[249] = 10'h35c;
        mem[250] = 10'h328;
        mem[251] = 10'h1eb;
        mem[252] = 10'h2b5;
        mem[253] = 10'h366;
        mem[254] = 10'h3f6;
        mem[255] = 10'h0bb;
        mem[256] = 10'h386;
        mem[257] = 10'h39c;
        mem[258] = 10'h3e2;
        mem[259] = 10'h1b2;
        mem[260] = 10'h0ce;
        mem[261] = 10'h21d;
        mem[262] = 10'h2ae;
        mem[263] = 10'h294;
        mem[264] = 10'h21f;
        mem[265] = 10'h1f3;
        mem[266] = 10'h1b7;
        mem[267] = 10'h313;
        mem[268] = 10'h166;
        mem[269] = 10'h3df;
        mem[270] = 10'h024;
        mem[271] = 10'h378;
        mem[272] = 10'h07e;
        mem[273] = 10'h2b9;
        mem[274] = 10'h29c;
        mem[275] = 10'h064;
        mem[276] = 10'h16b;
        mem[277] = 10'h2d6;
        mem[278] = 10'h309;
        mem[279] = 10'h11c;
        mem[280] = 10'h187;
        mem[281] = 10'h076;
        mem[282] = 10'h0be;
        mem[283] = 10'h36e;
        mem[284] = 10'h0db;
        mem[285] = 10'h165;
        mem[286] = 10'h19e;
        mem[287] = 10'h06c;
        mem[288] = 10'h39d;
        mem[289] = 10'h2fd;
        mem[290] = 10'h229;
        mem[291] = 10'h213;
        mem[292] = 10'h3ce;
        mem[293] = 10'h0ef;
        mem[294] = 10'h252;
        mem[295] = 10'h293;
        mem[296] = 10'h344;
        mem[297] = 10'h345;
        mem[298] = 10'h33a;
        mem[299] = 10'h15c;
        mem[300] = 10'h2f3;
        mem[301] = 10'h29a;
        mem[302] = 10'h116;
        mem[303] = 10'h1c1;
        mem[304] = 10'h095;
        mem[305] = 10'h261;
        mem[306] = 10'h1cc;
        mem[307] = 10'h2f4;
        mem[308] = 10'h0f7;
        mem[309] = 10'h0ff;
        mem[310] = 10'h1e5;
        mem[311] = 10'h23c;
        mem[312] = 10'h04f;
        mem[313] = 10'h283;
        mem[314] = 10'h15e;
        mem[315] = 10'h170;
        mem[316] = 10'h31a;
        mem[317] = 10'h2ca;
        mem[318] = 10'h2dc;
        mem[319] = 10'h2ad;
        mem[320] = 10'h1db;
        mem[321] = 10'h3ef;
        mem[322] = 10'h049;
        mem[323] = 10'h1a2;
        mem[324] = 10'h022;
        mem[325] = 10'h2ed;
        mem[326] = 10'h2ce;
        mem[327] = 10'h1fc;
        mem[328] = 10'h114;
        mem[329] = 10'h25f;
        mem[330] = 10'h2f0;
        mem[331] = 10'h195;
        mem[332] = 10'h330;
        mem[333] = 10'h3b6;
        mem[334] = 10'h07f;
        mem[335] = 10'h127;
        mem[336] = 10'h2e7;
        mem[337] = 10'h2f6;
        mem[338] = 10'h08e;
        mem[339] = 10'h398;
        mem[340] = 10'h227;
        mem[341] = 10'h3d0;
        mem[342] = 10'h0a5;
        mem[343] = 10'h1ec;
        mem[344] = 10'h092;
        mem[345] = 10'h1b9;
        mem[346] = 10'h007;
        mem[347] = 10'h38c;
        mem[348] = 10'h11d;
        mem[349] = 10'h03b;
        mem[350] = 10'h250;
        mem[351] = 10'h242;
        mem[352] = 10'h239;
        mem[353] = 10'h217;
        mem[354] = 10'h290;
        mem[355] = 10'h082;
        mem[356] = 10'h13c;
        mem[357] = 10'h123;
        mem[358] = 10'h28a;
        mem[359] = 10'h3e9;
        mem[360] = 10'h19f;
        mem[361] = 10'h35f;
        mem[362] = 10'h10f;
        mem[363] = 10'h09f;
        mem[364] = 10'h21c;
        mem[365] = 10'h3b3;
        mem[366] = 10'h373;
        mem[367] = 10'h385;
        mem[368] = 10'h1c0;
        mem[369] = 10'h380;
        mem[370] = 10'h140;
        mem[371] = 10'h21e;
        mem[372] = 10'h37a;
        mem[373] = 10'h120;
        mem[374] = 10'h1d5;
        mem[375] = 10'h375;
        mem[376] = 10'h14e;
        mem[377] = 10'h1de;
        mem[378] = 10'h13e;
        mem[379] = 10'h107;
        mem[380] = 10'h334;
        mem[381] = 10'h2f9;
        mem[382] = 10'h265;
        mem[383] = 10'h355;
        mem[384] = 10'h37c;
        mem[385] = 10'h01f;
        mem[386] = 10'h12d;
        mem[387] = 10'h01a;
        mem[388] = 10'h0a9;
        mem[389] = 10'h152;
        mem[390] = 10'h142;
        mem[391] = 10'h3dc;
        mem[392] = 10'h047;
        mem[393] = 10'h368;
        mem[394] = 10'h35b;
        mem[395] = 10'h230;
        mem[396] = 10'h33f;
        mem[397] = 10'h12f;
        mem[398] = 10'h108;
        mem[399] = 10'h002;
        mem[400] = 10'h2b7;
        mem[401] = 10'h26f;
        mem[402] = 10'h2bf;
        mem[403] = 10'h255;
        mem[404] = 10'h3ab;
        mem[405] = 10'h251;
        mem[406] = 10'h2cb;
        mem[407] = 10'h2fb;
        mem[408] = 10'h383;
        mem[409] = 10'h129;
        mem[410] = 10'h15b;
        mem[411] = 10'h3d4;
        mem[412] = 10'h102;
        mem[413] = 10'h01e;
        mem[414] = 10'h0e3;
        mem[415] = 10'h0a4;
        mem[416] = 10'h397;
        mem[417] = 10'h2c7;
        mem[418] = 10'h006;
        mem[419] = 10'h21b;
        mem[420] = 10'h22b;
        mem[421] = 10'h1df;
        mem[422] = 10'h22c;
        mem[423] = 10'h25d;
        mem[424] = 10'h238;
        mem[425] = 10'h2a3;
        mem[426] = 10'h2a0;
        mem[427] = 10'h138;
        mem[428] = 10'h192;
        mem[429] = 10'h15a;
        mem[430] = 10'h391;
        mem[431] = 10'h069;
        mem[432] = 10'h3e0;
        mem[433] = 10'h012;
        mem[434] = 10'h0b5;
        mem[435] = 10'h350;
        mem[436] = 10'h266;
        mem[437] = 10'h035;
        mem[438] = 10'h27c;
        mem[439] = 10'h0cb;
        mem[440] = 10'h008;
        mem[441] = 10'h38a;
        mem[442] = 10'h0cd;
        mem[443] = 10'h0fc;
        mem[444] = 10'h3d3;
        mem[445] = 10'h079;
        mem[446] = 10'h3ec;
        mem[447] = 10'h148;
        mem[448] = 10'h2c6;
        mem[449] = 10'h324;
        mem[450] = 10'h122;
        mem[451] = 10'h11f;
        mem[452] = 10'h161;
        mem[453] = 10'h202;
        mem[454] = 10'h3db;
        mem[455] = 10'h2e5;
        mem[456] = 10'h0ae;
        mem[457] = 10'h12b;
        mem[458] = 10'h2c8;
        mem[459] = 10'h2e4;
        mem[460] = 10'h263;
        mem[461] = 10'h2b0;
        mem[462] = 10'h1cb;
        mem[463] = 10'h0f5;
        mem[464] = 10'h30b;
        mem[465] = 10'h09e;
        mem[466] = 10'h284;
        mem[467] = 10'h3a2;
        mem[468] = 10'h00b;
        mem[469] = 10'h030;
        mem[470] = 10'h05b;
        mem[471] = 10'h091;
        mem[472] = 10'h302;
        mem[473] = 10'h2d4;
        mem[474] = 10'h236;
        mem[475] = 10'h3cb;
        mem[476] = 10'h316;
        mem[477] = 10'h16f;
        mem[478] = 10'h098;
        mem[479] = 10'h02a;
        mem[480] = 10'h077;
        mem[481] = 10'h3b5;
        mem[482] = 10'h0c5;
        mem[483] = 10'h0cf;
        mem[484] = 10'h167;
        mem[485] = 10'h3bc;
        mem[486] = 10'h057;
        mem[487] = 10'h04a;
        mem[488] = 10'h0b9;
        mem[489] = 10'h287;
        mem[490] = 10'h10b;
        mem[491] = 10'h1bb;
        mem[492] = 10'h2df;
        mem[493] = 10'h015;
        mem[494] = 10'h0d2;
        mem[495] = 10'h0d3;
        mem[496] = 10'h03d;
        mem[497] = 10'h221;
        mem[498] = 10'h1c6;
        mem[499] = 10'h3c8;
        mem[500] = 10'h228;
        mem[501] = 10'h342;
        mem[502] = 10'h353;
        mem[503] = 10'h2c3;
        mem[504] = 10'h315;
        mem[505] = 10'h370;
        mem[506] = 10'h0c2;
        mem[507] = 10'h0f6;
        mem[508] = 10'h3c9;
        mem[509] = 10'h20c;
        mem[510] = 10'h174;
        mem[511] = 10'h1d4;
        mem[512] = 10'h3e3;
        mem[513] = 10'h23e;
        mem[514] = 10'h132;
        mem[515] = 10'h3f3;
        mem[516] = 10'h2a5;
        mem[517] = 10'h3a5;
        mem[518] = 10'h26b;
        mem[519] = 10'h15d;
        mem[520] = 10'h089;
        mem[521] = 10'h29d;
        mem[522] = 10'h393;
        mem[523] = 10'h3ee;
        mem[524] = 10'h3e6;
        mem[525] = 10'h27d;
        mem[526] = 10'h1e0;
        mem[527] = 10'h0d5;
        mem[528] = 10'h308;
        mem[529] = 10'h3c2;
        mem[530] = 10'h097;
        mem[531] = 10'h319;
        mem[532] = 10'h042;
        mem[533] = 10'h08d;
        mem[534] = 10'h1fb;
        mem[535] = 10'h033;
        mem[536] = 10'h3f8;
        mem[537] = 10'h292;
        mem[538] = 10'h17d;
        mem[539] = 10'h323;
        mem[540] = 10'h341;
        mem[541] = 10'h39b;
        mem[542] = 10'h00c;
        mem[543] = 10'h399;
        mem[544] = 10'h080;
        mem[545] = 10'h1ef;
        mem[546] = 10'h0df;
        mem[547] = 10'h367;
        mem[548] = 10'h295;
        mem[549] = 10'h018;
        mem[550] = 10'h23b;
        mem[551] = 10'h193;
        mem[552] = 10'h20d;
        mem[553] = 10'h131;
        mem[554] = 10'h0d1;
        mem[555] = 10'h037;
        mem[556] = 10'h155;
        mem[557] = 10'h000;
        mem[558] = 10'h338;
        mem[559] = 10'h32f;
        mem[560] = 10'h093;
        mem[561] = 10'h065;
        mem[562] = 10'h0c9;
        mem[563] = 10'h365;
        mem[564] = 10'h320;
        mem[565] = 10'h09a;
        mem[566] = 10'h28b;
        mem[567] = 10'h34a;
        mem[568] = 10'h26e;
        mem[569] = 10'h11e;
        mem[570] = 10'h3a0;
        mem[571] = 10'h207;
        mem[572] = 10'h05d;
        mem[573] = 10'h2fc;
        mem[574] = 10'h0aa;
        mem[575] = 10'h210;
        mem[576] = 10'h1b3;
        mem[577] = 10'h2ac;
        mem[578] = 10'h31b;
        mem[579] = 10'h0ed;
        mem[580] = 10'h0fa;
        mem[581] = 10'h13d;
        mem[582] = 10'h02f;
        mem[583] = 10'h347;
        mem[584] = 10'h201;
        mem[585] = 10'h04e;
        mem[586] = 10'h32e;
        mem[587] = 10'h02d;
        mem[588] = 10'h073;
        mem[589] = 10'h0a7;
        mem[590] = 10'h07d;
        mem[591] = 10'h040;
        mem[592] = 10'h282;
        mem[593] = 10'h214;
        mem[594] = 10'h1f8;
        mem[595] = 10'h2a8;
        mem[596] = 10'h310;
        mem[597] = 10'h211;
        mem[598] = 10'h26d;
        mem[599] = 10'h24f;
        mem[600] = 10'h2bb;
        mem[601] = 10'h178;
        mem[602] = 10'h262;
        mem[603] = 10'h392;
        mem[604] = 10'h29f;
        mem[605] = 10'h357;
        mem[606] = 10'h276;
        mem[607] = 10'h33b;
        mem[608] = 10'h08f;
        mem[609] = 10'h130;
        mem[610] = 10'h1dc;
        mem[611] = 10'h0c7;
        mem[612] = 10'h3a4;
        mem[613] = 10'h23d;
        mem[614] = 10'h3af;
        mem[615] = 10'h2c0;
        mem[616] = 10'h173;
        mem[617] = 10'h1f0;
        mem[618] = 10'h1aa;
        mem[619] = 10'h33c;
        mem[620] = 10'h1a1;
        mem[621] = 10'h2af;
        mem[622] = 10'h0a1;
        mem[623] = 10'h24e;
        mem[624] = 10'h271;
        mem[625] = 10'h2e3;
        mem[626] = 10'h0fe;
        mem[627] = 10'h1d1;
        mem[628] = 10'h181;
        mem[629] = 10'h22f;
        mem[630] = 10'h14d;
        mem[631] = 10'h197;
        mem[632] = 10'h094;
        mem[633] = 10'h02b;
        mem[634] = 10'h1f4;
        mem[635] = 10'h00e;
        mem[636] = 10'h34e;
        mem[637] = 10'h1a6;
        mem[638] = 10'h3d8;
        mem[639] = 10'h1be;
        mem[640] = 10'h10d;
        mem[641] = 10'h390;
        mem[642] = 10'h081;
        mem[643] = 10'h24c;
        mem[644] = 10'h2a6;
        mem[645] = 10'h2d9;
        mem[646] = 10'h289;
        mem[647] = 10'h31c;
        mem[648] = 10'h3a1;
        mem[649] = 10'h067;
        mem[650] = 10'h1af;
        mem[651] = 10'h013;
        mem[652] = 10'h1da;
        mem[653] = 10'h0dc;
        mem[654] = 10'h2cc;
        mem[655] = 10'h16d;
        mem[656] = 10'h032;
        mem[657] = 10'h3b8;
        mem[658] = 10'h021;
        mem[659] = 10'h09c;
        mem[660] = 10'h189;
        mem[661] = 10'h2fe;
        mem[662] = 10'h2d1;
        mem[663] = 10'h17b;
        mem[664] = 10'h3ff;
        mem[665] = 10'h2c9;
        mem[666] = 10'h0b0;
        mem[667] = 10'h16e;
        mem[668] = 10'h31d;
        mem[669] = 10'h07b;
        mem[670] = 10'h34c;
        mem[671] = 10'h200;
        mem[672] = 10'h25b;
        mem[673] = 10'h3a7;
        mem[674] = 10'h06e;
        mem[675] = 10'h044;
        mem[676] = 10'h03e;
        mem[677] = 10'h01d;
        mem[678] = 10'h306;
        mem[679] = 10'h269;
        mem[680] = 10'h3b0;
        mem[681] = 10'h185;
        mem[682] = 10'h395;
        mem[683] = 10'h025;
        mem[684] = 10'h216;
        mem[685] = 10'h0f0;
        mem[686] = 10'h1f6;
        mem[687] = 10'h18c;
        mem[688] = 10'h02e;
        mem[689] = 10'h128;
        mem[690] = 10'h3be;
        mem[691] = 10'h068;
        mem[692] = 10'h001;
        mem[693] = 10'h30a;
        mem[694] = 10'h17c;
        mem[695] = 10'h0bf;
        mem[696] = 10'h28f;
        mem[697] = 10'h050;
        mem[698] = 10'h052;
        mem[699] = 10'h0a2;
        mem[700] = 10'h009;
        mem[701] = 10'h3dd;
        mem[702] = 10'h088;
        mem[703] = 10'h14a;
        mem[704] = 10'h005;
        mem[705] = 10'h00a;
        mem[706] = 10'h0bd;
        mem[707] = 10'h0da;
        mem[708] = 10'h34b;
        mem[709] = 10'h332;
        mem[710] = 10'h0ee;
        mem[711] = 10'h19b;
        mem[712] = 10'h0e7;
        mem[713] = 10'h329;
        mem[714] = 10'h225;
        mem[715] = 10'h110;
        mem[716] = 10'h360;
        mem[717] = 10'h18b;
        mem[718] = 10'h2dd;
        mem[719] = 10'h3d9;
        mem[720] = 10'h321;
        mem[721] = 10'h3bd;
        mem[722] = 10'h0c0;
        mem[723] = 10'h3de;
        mem[724] = 10'h387;
        mem[725] = 10'h325;
        mem[726] = 10'h126;
        mem[727] = 10'h0b4;
        mem[728] = 10'h1b8;
        mem[729] = 10'h3f4;
        mem[730] = 10'h0cc;
        mem[731] = 10'h2ea;
        mem[732] = 10'h233;
        mem[733] = 10'h298;
        mem[734] = 10'h291;
        mem[735] = 10'h059;
        mem[736] = 10'h0d8;
        mem[737] = 10'h1ac;
        mem[738] = 10'h124;
        mem[739] = 10'h30d;
        mem[740] = 10'h0bc;
        mem[741] = 10'h053;
        mem[742] = 10'h247;
        mem[743] = 10'h2c1;
        mem[744] = 10'h249;
        mem[745] = 10'h384;
        mem[746] = 10'h0e6;
        mem[747] = 10'h352;
        mem[748] = 10'h37f;
        mem[749] = 10'h0f3;
        mem[750] = 10'h074;
        mem[751] = 10'h1fd;
        mem[752] = 10'h218;
        mem[753] = 10'h281;
        mem[754] = 10'h186;
        mem[755] = 10'h1cf;
        mem[756] = 10'h2cf;
        mem[757] = 10'h070;
        mem[758] = 10'h18d;
        mem[759] = 10'h172;
        mem[760] = 10'h096;
        mem[761] = 10'h06f;
        mem[762] = 10'h3eb;
        mem[763] = 10'h38e;
        mem[764] = 10'h36f;
        mem[765] = 10'h169;
        mem[766] = 10'h300;
        mem[767] = 10'h099;
        mem[768] = 10'h1d3;
        mem[769] = 10'h1c4;
        mem[770] = 10'h0b2;
        mem[771] = 10'h3fc;
        mem[772] = 10'h235;
        mem[773] = 10'h3e1;
        mem[774] = 10'h3c5;
        mem[775] = 10'h336;
        mem[776] = 10'h27e;
        mem[777] = 10'h0c1;
        mem[778] = 10'h13b;
        mem[779] = 10'h149;
        mem[780] = 10'h1ee;
        mem[781] = 10'h3a8;
        mem[782] = 10'h19a;
        mem[783] = 10'h299;
        mem[784] = 10'h153;
        mem[785] = 10'h144;
        mem[786] = 10'h121;
        mem[787] = 10'h1d2;
        mem[788] = 10'h27f;
        mem[789] = 10'h2ef;
        mem[790] = 10'h3fb;
        mem[791] = 10'h190;
        mem[792] = 10'h27b;
        mem[793] = 10'h2b2;
        mem[794] = 10'h3c6;
        mem[795] = 10'h30e;
        mem[796] = 10'h35a;
        mem[797] = 10'h1fa;
        mem[798] = 10'h246;
        mem[799] = 10'h3c3;
        mem[800] = 10'h1e2;
        mem[801] = 10'h286;
        mem[802] = 10'h272;
        mem[803] = 10'h118;
        mem[804] = 10'h25c;
        mem[805] = 10'h396;
        mem[806] = 10'h35d;
        mem[807] = 10'h0e5;
        mem[808] = 10'h06d;
        mem[809] = 10'h22a;
        mem[810] = 10'h29e;
        mem[811] = 10'h0f2;
        mem[812] = 10'h0d0;
        mem[813] = 10'h268;
        mem[814] = 10'h046;
        mem[815] = 10'h196;
        mem[816] = 10'h296;
        mem[817] = 10'h163;
        mem[818] = 10'h220;
        mem[819] = 10'h179;
        mem[820] = 10'h1c2;
        mem[821] = 10'h05f;
        mem[822] = 10'h3f5;
        mem[823] = 10'h24d;
        mem[824] = 10'h0d6;
        mem[825] = 10'h084;
        mem[826] = 10'h04b;
        mem[827] = 10'h318;
        mem[828] = 10'h326;
        mem[829] = 10'h2b6;
        mem[830] = 10'h17a;
        mem[831] = 10'h285;
        mem[832] = 10'h369;
        mem[833] = 10'h376;
        mem[834] = 10'h020;
        mem[835] = 10'h25e;
        mem[836] = 10'h1a8;
        mem[837] = 10'h0d4;
        mem[838] = 10'h0e8;
        mem[839] = 10'h1ab;
        mem[840] = 10'h3a9;
        mem[841] = 10'h20a;
        mem[842] = 10'h38f;
        mem[843] = 10'h23a;
        mem[844] = 10'h206;
        mem[845] = 10'h058;
        mem[846] = 10'h0b7;
        mem[847] = 10'h1d9;
        mem[848] = 10'h24b;
        mem[849] = 10'h2a1;
        mem[850] = 10'h3d2;
        mem[851] = 10'h231;
        mem[852] = 10'h223;
        mem[853] = 10'h297;
        mem[854] = 10'h32b;
        mem[855] = 10'h257;
        mem[856] = 10'h16c;
        mem[857] = 10'h2a7;
        mem[858] = 10'h0b6;
        mem[859] = 10'h1ca;
        mem[860] = 10'h1e4;
        mem[861] = 10'h0c6;
        mem[862] = 10'h2f7;
        mem[863] = 10'h09d;
        mem[864] = 10'h32d;
        mem[865] = 10'h019;
        mem[866] = 10'h1f1;
        mem[867] = 10'h331;
        mem[868] = 10'h085;
        mem[869] = 10'h1fe;
        mem[870] = 10'h164;
        mem[871] = 10'h3c4;
        mem[872] = 10'h1e8;
        mem[873] = 10'h156;
        mem[874] = 10'h1ed;
        mem[875] = 10'h0eb;
        mem[876] = 10'h3f2;
        mem[877] = 10'h0b3;
        mem[878] = 10'h101;
        mem[879] = 10'h2ab;
        mem[880] = 10'h3d5;
        mem[881] = 10'h10c;
        mem[882] = 10'h1d0;
        mem[883] = 10'h1c8;
        mem[884] = 10'h3d7;
        mem[885] = 10'h348;
        mem[886] = 10'h22e;
        mem[887] = 10'h18a;
        mem[888] = 10'h20f;
        mem[889] = 10'h0fd;
        mem[890] = 10'h224;
        mem[891] = 10'h1c5;
        mem[892] = 10'h056;
        mem[893] = 10'h38b;
        mem[894] = 10'h205;
        mem[895] = 10'h2f1;
        mem[896] = 10'h2e0;
        mem[897] = 10'h00d;
        mem[898] = 10'h374;
        mem[899] = 10'h04d;
        mem[900] = 10'h3ba;
        mem[901] = 10'h1bc;
        mem[902] = 10'h3e8;
        mem[903] = 10'h0c3;
        mem[904] = 10'h111;
        mem[905] = 10'h3e4;
        mem[906] = 10'h258;
        mem[907] = 10'h394;
        mem[908] = 10'h105;
        mem[909] = 10'h2a9;
        mem[910] = 10'h232;
        mem[911] = 10'h25a;
        mem[912] = 10'h038;
        mem[913] = 10'h3ae;
        mem[914] = 10'h3fa;
        mem[915] = 10'h01c;
        mem[916] = 10'h1a0;
        mem[917] = 10'h0e9;
        mem[918] = 10'h3ea;
        mem[919] = 10'h2eb;
        mem[920] = 10'h028;
        mem[921] = 10'h026;
        mem[922] = 10'h3e5;
        mem[923] = 10'h260;
        mem[924] = 10'h18f;
        mem[925] = 10'h175;
        mem[926] = 10'h075;
        mem[927] = 10'h3b7;
        mem[928] = 10'h1e1;
        mem[929] = 10'h100;
        mem[930] = 10'h362;
        mem[931] = 10'h3ad;
        mem[932] = 10'h22d;
        mem[933] = 10'h2f2;
        mem[934] = 10'h066;
        mem[935] = 10'h311;
        mem[936] = 10'h1b6;
        mem[937] = 10'h3fd;
        mem[938] = 10'h183;
        mem[939] = 10'h03f;
        mem[940] = 10'h06a;
        mem[941] = 10'h2fa;
        mem[942] = 10'h16a;
        mem[943] = 10'h1f2;
        mem[944] = 10'h1e9;
        mem[945] = 10'h1a5;
        mem[946] = 10'h11b;
        mem[947] = 10'h3b1;
        mem[948] = 10'h3f9;
        mem[949] = 10'h35e;
        mem[950] = 10'h273;
        mem[951] = 10'h0d9;
        mem[952] = 10'h1e7;
        mem[953] = 10'h145;
        mem[954] = 10'h275;
        mem[955] = 10'h3ac;
        mem[956] = 10'h2e1;
        mem[957] = 10'h1ad;
        mem[958] = 10'h358;
        mem[959] = 10'h051;
        mem[960] = 10'h2e8;
        mem[961] = 10'h2b4;
        mem[962] = 10'h07a;
        mem[963] = 10'h188;
        mem[964] = 10'h3cc;
        mem[965] = 10'h055;
        mem[966] = 10'h176;
        mem[967] = 10'h0ca;
        mem[968] = 10'h2d7;
        mem[969] = 10'h3f1;
        mem[970] = 10'h199;
        mem[971] = 10'h2ff;
        mem[972] = 10'h0e4;
        mem[973] = 10'h12e;
        mem[974] = 10'h003;
        mem[975] = 10'h05e;
        mem[976] = 10'h1e6;
        mem[977] = 10'h2aa;
        mem[978] = 10'h3f0;
        mem[979] = 10'h031;
        mem[980] = 10'h361;
        mem[981] = 10'h1d6;
        mem[982] = 10'h04c;
        mem[983] = 10'h30f;
        mem[984] = 10'h377;
        mem[985] = 10'h119;
        mem[986] = 10'h240;
        mem[987] = 10'h1cd;
        mem[988] = 10'h1ea;
        mem[989] = 10'h029;
        mem[990] = 10'h24a;
        mem[991] = 10'h00f;
        mem[992] = 10'h115;
        mem[993] = 10'h209;
        mem[994] = 10'h215;
        mem[995] = 10'h2d3;
        mem[996] = 10'h0f9;
        mem[997] = 10'h054;
        mem[998] = 10'h13a;
        mem[999] = 10'h379;
        mem[1000] = 10'h3aa;
        mem[1001] = 10'h17f;
        mem[1002] = 10'h3da;
        mem[1003] = 10'h087;
        mem[1004] = 10'h31f;
        mem[1005] = 10'h1b4;
        mem[1006] = 10'h0a6;
        mem[1007] = 10'h14b;
        mem[1008] = 10'h34d;
        mem[1009] = 10'h314;
        mem[1010] = 10'h0ad;
        mem[1011] = 10'h359;
        mem[1012] = 10'h1d7;
        mem[1013] = 10'h33e;
        mem[1014] = 10'h1f7;
        mem[1015] = 10'h1dd;
        mem[1016] = 10'h1ba;
        mem[1017] = 10'h307;
        mem[1018] = 10'h0b1;
        mem[1019] = 10'h1bf;
        mem[1020] = 10'h08b;
        mem[1021] = 10'h0c4;
        mem[1022] = 10'h182;
        mem[1023] = 10'h13f;
    end
endmodule

module odo_apply_sboxes(clk, in, out);
    input clk;
    input [639:0] in;
    output [639:0] out;
    odo_sbox_small0 sbox0inst(clk, in[5:0], out[5:0]);
    odo_sbox_small1 sbox1inst(clk, in[21:16], out[21:16]);
    odo_sbox_large0 sbox2inst(clk, in[15:6], in[31:22], out[15:6], out[31:22]);
    odo_sbox_small2 sbox3inst(clk, in[37:32], out[37:32]);
    odo_sbox_small3 sbox4inst(clk, in[53:48], out[53:48]);
    odo_sbox_large0 sbox5inst(clk, in[47:38], in[63:54], out[47:38], out[63:54]);
    odo_sbox_small4 sbox6inst(clk, in[69:64], out[69:64]);
    odo_sbox_small5 sbox7inst(clk, in[85:80], out[85:80]);
    odo_sbox_large1 sbox8inst(clk, in[79:70], in[95:86], out[79:70], out[95:86]);
    odo_sbox_small6 sbox9inst(clk, in[101:96], out[101:96]);
    odo_sbox_small7 sbox10inst(clk, in[117:112], out[117:112]);
    odo_sbox_large1 sbox11inst(clk, in[111:102], in[127:118], out[111:102], out[127:118]);
    odo_sbox_small8 sbox12inst(clk, in[133:128], out[133:128]);
    odo_sbox_small9 sbox13inst(clk, in[149:144], out[149:144]);
    odo_sbox_large2 sbox14inst(clk, in[143:134], in[159:150], out[143:134], out[159:150]);
    odo_sbox_small10 sbox15inst(clk, in[165:160], out[165:160]);
    odo_sbox_small11 sbox16inst(clk, in[181:176], out[181:176]);
    odo_sbox_large2 sbox17inst(clk, in[175:166], in[191:182], out[175:166], out[191:182]);
    odo_sbox_small12 sbox18inst(clk, in[197:192], out[197:192]);
    odo_sbox_small13 sbox19inst(clk, in[213:208], out[213:208]);
    odo_sbox_large3 sbox20inst(clk, in[207:198], in[223:214], out[207:198], out[223:214]);
    odo_sbox_small14 sbox21inst(clk, in[229:224], out[229:224]);
    odo_sbox_small15 sbox22inst(clk, in[245:240], out[245:240]);
    odo_sbox_large3 sbox23inst(clk, in[239:230], in[255:246], out[239:230], out[255:246]);
    odo_sbox_small16 sbox24inst(clk, in[261:256], out[261:256]);
    odo_sbox_small17 sbox25inst(clk, in[277:272], out[277:272]);
    odo_sbox_large4 sbox26inst(clk, in[271:262], in[287:278], out[271:262], out[287:278]);
    odo_sbox_small18 sbox27inst(clk, in[293:288], out[293:288]);
    odo_sbox_small19 sbox28inst(clk, in[309:304], out[309:304]);
    odo_sbox_large4 sbox29inst(clk, in[303:294], in[319:310], out[303:294], out[319:310]);
    odo_sbox_small20 sbox30inst(clk, in[325:320], out[325:320]);
    odo_sbox_small21 sbox31inst(clk, in[341:336], out[341:336]);
    odo_sbox_large5 sbox32inst(clk, in[335:326], in[351:342], out[335:326], out[351:342]);
    odo_sbox_small22 sbox33inst(clk, in[357:352], out[357:352]);
    odo_sbox_small23 sbox34inst(clk, in[373:368], out[373:368]);
    odo_sbox_large5 sbox35inst(clk, in[367:358], in[383:374], out[367:358], out[383:374]);
    odo_sbox_small24 sbox36inst(clk, in[389:384], out[389:384]);
    odo_sbox_small25 sbox37inst(clk, in[405:400], out[405:400]);
    odo_sbox_large6 sbox38inst(clk, in[399:390], in[415:406], out[399:390], out[415:406]);
    odo_sbox_small26 sbox39inst(clk, in[421:416], out[421:416]);
    odo_sbox_small27 sbox40inst(clk, in[437:432], out[437:432]);
    odo_sbox_large6 sbox41inst(clk, in[431:422], in[447:438], out[431:422], out[447:438]);
    odo_sbox_small28 sbox42inst(clk, in[453:448], out[453:448]);
    odo_sbox_small29 sbox43inst(clk, in[469:464], out[469:464]);
    odo_sbox_large7 sbox44inst(clk, in[463:454], in[479:470], out[463:454], out[479:470]);
    odo_sbox_small30 sbox45inst(clk, in[485:480], out[485:480]);
    odo_sbox_small31 sbox46inst(clk, in[501:496], out[501:496]);
    odo_sbox_large7 sbox47inst(clk, in[495:486], in[511:502], out[495:486], out[511:502]);
    odo_sbox_small32 sbox48inst(clk, in[517:512], out[517:512]);
    odo_sbox_small33 sbox49inst(clk, in[533:528], out[533:528]);
    odo_sbox_large8 sbox50inst(clk, in[527:518], in[543:534], out[527:518], out[543:534]);
    odo_sbox_small34 sbox51inst(clk, in[549:544], out[549:544]);
    odo_sbox_small35 sbox52inst(clk, in[565:560], out[565:560]);
    odo_sbox_large8 sbox53inst(clk, in[559:550], in[575:566], out[559:550], out[575:566]);
    odo_sbox_small36 sbox54inst(clk, in[581:576], out[581:576]);
    odo_sbox_small37 sbox55inst(clk, in[597:592], out[597:592]);
    odo_sbox_large9 sbox56inst(clk, in[591:582], in[607:598], out[591:582], out[607:598]);
    odo_sbox_small38 sbox57inst(clk, in[613:608], out[613:608]);
    odo_sbox_small39 sbox58inst(clk, in[629:624], out[629:624]);
    odo_sbox_large9 sbox59inst(clk, in[623:614], in[639:630], out[623:614], out[639:630]);
endmodule

module odo_apply_pbox0(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[444] = in[0];
    assign out[83] = in[1];
    assign out[324] = in[2];
    assign out[350] = in[3];
    assign out[21] = in[4];
    assign out[405] = in[5];
    assign out[66] = in[6];
    assign out[265] = in[7];
    assign out[496] = in[8];
    assign out[208] = in[9];
    assign out[228] = in[10];
    assign out[540] = in[11];
    assign out[72] = in[12];
    assign out[393] = in[13];
    assign out[213] = in[14];
    assign out[32] = in[15];
    assign out[480] = in[16];
    assign out[196] = in[17];
    assign out[14] = in[18];
    assign out[173] = in[19];
    assign out[400] = in[20];
    assign out[343] = in[21];
    assign out[157] = in[22];
    assign out[410] = in[23];
    assign out[60] = in[24];
    assign out[489] = in[25];
    assign out[201] = in[26];
    assign out[414] = in[27];
    assign out[452] = in[28];
    assign out[327] = in[29];
    assign out[519] = in[30];
    assign out[185] = in[31];
    assign out[633] = in[32];
    assign out[11] = in[33];
    assign out[635] = in[34];
    assign out[539] = in[35];
    assign out[613] = in[36];
    assign out[352] = in[37];
    assign out[55] = in[38];
    assign out[57] = in[39];
    assign out[234] = in[40];
    assign out[618] = in[41];
    assign out[466] = in[42];
    assign out[171] = in[43];
    assign out[499] = in[44];
    assign out[279] = in[45];
    assign out[341] = in[46];
    assign out[19] = in[47];
    assign out[585] = in[48];
    assign out[500] = in[49];
    assign out[514] = in[50];
    assign out[29] = in[51];
    assign out[347] = in[52];
    assign out[582] = in[53];
    assign out[144] = in[54];
    assign out[435] = in[55];
    assign out[167] = in[56];
    assign out[236] = in[57];
    assign out[611] = in[58];
    assign out[48] = in[59];
    assign out[131] = in[60];
    assign out[614] = in[61];
    assign out[442] = in[62];
    assign out[527] = in[63];
    assign out[295] = in[64];
    assign out[456] = in[65];
    assign out[300] = in[66];
    assign out[221] = in[67];
    assign out[203] = in[68];
    assign out[597] = in[69];
    assign out[583] = in[70];
    assign out[639] = in[71];
    assign out[202] = in[72];
    assign out[562] = in[73];
    assign out[397] = in[74];
    assign out[333] = in[75];
    assign out[541] = in[76];
    assign out[360] = in[77];
    assign out[615] = in[78];
    assign out[632] = in[79];
    assign out[584] = in[80];
    assign out[235] = in[81];
    assign out[571] = in[82];
    assign out[37] = in[83];
    assign out[56] = in[84];
    assign out[38] = in[85];
    assign out[337] = in[86];
    assign out[624] = in[87];
    assign out[339] = in[88];
    assign out[224] = in[89];
    assign out[406] = in[90];
    assign out[482] = in[91];
    assign out[24] = in[92];
    assign out[542] = in[93];
    assign out[598] = in[94];
    assign out[91] = in[95];
    assign out[521] = in[96];
    assign out[561] = in[97];
    assign out[6] = in[98];
    assign out[117] = in[99];
    assign out[604] = in[100];
    assign out[332] = in[101];
    assign out[321] = in[102];
    assign out[430] = in[103];
    assign out[335] = in[104];
    assign out[101] = in[105];
    assign out[595] = in[106];
    assign out[572] = in[107];
    assign out[637] = in[108];
    assign out[367] = in[109];
    assign out[99] = in[110];
    assign out[177] = in[111];
    assign out[267] = in[112];
    assign out[429] = in[113];
    assign out[281] = in[114];
    assign out[431] = in[115];
    assign out[187] = in[116];
    assign out[181] = in[117];
    assign out[90] = in[118];
    assign out[520] = in[119];
    assign out[447] = in[120];
    assign out[251] = in[121];
    assign out[531] = in[122];
    assign out[170] = in[123];
    assign out[451] = in[124];
    assign out[189] = in[125];
    assign out[104] = in[126];
    assign out[576] = in[127];
    assign out[315] = in[128];
    assign out[348] = in[129];
    assign out[535] = in[130];
    assign out[467] = in[131];
    assign out[404] = in[132];
    assign out[127] = in[133];
    assign out[555] = in[134];
    assign out[45] = in[135];
    assign out[0] = in[136];
    assign out[389] = in[137];
    assign out[293] = in[138];
    assign out[411] = in[139];
    assign out[70] = in[140];
    assign out[214] = in[141];
    assign out[458] = in[142];
    assign out[548] = in[143];
    assign out[209] = in[144];
    assign out[510] = in[145];
    assign out[269] = in[146];
    assign out[395] = in[147];
    assign out[355] = in[148];
    assign out[318] = in[149];
    assign out[319] = in[150];
    assign out[264] = in[151];
    assign out[155] = in[152];
    assign out[162] = in[153];
    assign out[490] = in[154];
    assign out[263] = in[155];
    assign out[468] = in[156];
    assign out[605] = in[157];
    assign out[459] = in[158];
    assign out[460] = in[159];
    assign out[601] = in[160];
    assign out[432] = in[161];
    assign out[434] = in[162];
    assign out[498] = in[163];
    assign out[210] = in[164];
    assign out[308] = in[165];
    assign out[373] = in[166];
    assign out[77] = in[167];
    assign out[153] = in[168];
    assign out[260] = in[169];
    assign out[553] = in[170];
    assign out[546] = in[171];
    assign out[506] = in[172];
    assign out[222] = in[173];
    assign out[241] = in[174];
    assign out[288] = in[175];
    assign out[284] = in[176];
    assign out[554] = in[177];
    assign out[365] = in[178];
    assign out[416] = in[179];
    assign out[231] = in[180];
    assign out[522] = in[181];
    assign out[523] = in[182];
    assign out[631] = in[183];
    assign out[525] = in[184];
    assign out[606] = in[185];
    assign out[363] = in[186];
    assign out[592] = in[187];
    assign out[394] = in[188];
    assign out[566] = in[189];
    assign out[54] = in[190];
    assign out[462] = in[191];
    assign out[137] = in[192];
    assign out[362] = in[193];
    assign out[569] = in[194];
    assign out[443] = in[195];
    assign out[557] = in[196];
    assign out[256] = in[197];
    assign out[303] = in[198];
    assign out[106] = in[199];
    assign out[407] = in[200];
    assign out[314] = in[201];
    assign out[139] = in[202];
    assign out[49] = in[203];
    assign out[388] = in[204];
    assign out[497] = in[205];
    assign out[215] = in[206];
    assign out[477] = in[207];
    assign out[565] = in[208];
    assign out[218] = in[209];
    assign out[379] = in[210];
    assign out[354] = in[211];
    assign out[151] = in[212];
    assign out[257] = in[213];
    assign out[124] = in[214];
    assign out[154] = in[215];
    assign out[422] = in[216];
    assign out[220] = in[217];
    assign out[262] = in[218];
    assign out[156] = in[219];
    assign out[165] = in[220];
    assign out[518] = in[221];
    assign out[204] = in[222];
    assign out[600] = in[223];
    assign out[629] = in[224];
    assign out[25] = in[225];
    assign out[147] = in[226];
    assign out[475] = in[227];
    assign out[351] = in[228];
    assign out[481] = in[229];
    assign out[418] = in[230];
    assign out[310] = in[231];
    assign out[438] = in[232];
    assign out[440] = in[233];
    assign out[80] = in[234];
    assign out[487] = in[235];
    assign out[280] = in[236];
    assign out[182] = in[237];
    assign out[445] = in[238];
    assign out[423] = in[239];
    assign out[345] = in[240];
    assign out[364] = in[241];
    assign out[42] = in[242];
    assign out[322] = in[243];
    assign out[46] = in[244];
    assign out[254] = in[245];
    assign out[453] = in[246];
    assign out[484] = in[247];
    assign out[193] = in[248];
    assign out[328] = in[249];
    assign out[591] = in[250];
    assign out[356] = in[251];
    assign out[504] = in[252];
    assign out[312] = in[253];
    assign out[172] = in[254];
    assign out[240] = in[255];
    assign out[479] = in[256];
    assign out[178] = in[257];
    assign out[586] = in[258];
    assign out[244] = in[259];
    assign out[574] = in[260];
    assign out[64] = in[261];
    assign out[616] = in[262];
    assign out[184] = in[263];
    assign out[494] = in[264];
    assign out[78] = in[265];
    assign out[105] = in[266];
    assign out[296] = in[267];
    assign out[369] = in[268];
    assign out[298] = in[269];
    assign out[270] = in[270];
    assign out[102] = in[271];
    assign out[103] = in[272];
    assign out[40] = in[273];
    assign out[533] = in[274];
    assign out[545] = in[275];
    assign out[43] = in[276];
    assign out[247] = in[277];
    assign out[538] = in[278];
    assign out[249] = in[279];
    assign out[426] = in[280];
    assign out[382] = in[281];
    assign out[121] = in[282];
    assign out[313] = in[283];
    assign out[304] = in[284];
    assign out[544] = in[285];
    assign out[39] = in[286];
    assign out[577] = in[287];
    assign out[552] = in[288];
    assign out[175] = in[289];
    assign out[383] = in[290];
    assign out[448] = in[291];
    assign out[252] = in[292];
    assign out[470] = in[293];
    assign out[622] = in[294];
    assign out[108] = in[295];
    assign out[71] = in[296];
    assign out[474] = in[297];
    assign out[508] = in[298];
    assign out[476] = in[299];
    assign out[344] = in[300];
    assign out[12] = in[301];
    assign out[41] = in[302];
    assign out[593] = in[303];
    assign out[461] = in[304];
    assign out[628] = in[305];
    assign out[399] = in[306];
    assign out[297] = in[307];
    assign out[75] = in[308];
    assign out[309] = in[309];
    assign out[412] = in[310];
    assign out[227] = in[311];
    assign out[226] = in[312];
    assign out[62] = in[313];
    assign out[3] = in[314];
    assign out[472] = in[315];
    assign out[168] = in[316];
    assign out[174] = in[317];
    assign out[239] = in[318];
    assign out[349] = in[319];
    assign out[31] = in[320];
    assign out[207] = in[321];
    assign out[134] = in[322];
    assign out[323] = in[323];
    assign out[530] = in[324];
    assign out[325] = in[325];
    assign out[292] = in[326];
    assign out[485] = in[327];
    assign out[588] = in[328];
    assign out[186] = in[329];
    assign out[526] = in[330];
    assign out[517] = in[331];
    assign out[81] = in[332];
    assign out[115] = in[333];
    assign out[116] = in[334];
    assign out[417] = in[335];
    assign out[502] = in[336];
    assign out[596] = in[337];
    assign out[23] = in[338];
    assign out[421] = in[339];
    assign out[122] = in[340];
    assign out[191] = in[341];
    assign out[488] = in[342];
    assign out[125] = in[343];
    assign out[501] = in[344];
    assign out[34] = in[345];
    assign out[35] = in[346];
    assign out[135] = in[347];
    assign out[507] = in[348];
    assign out[609] = in[349];
    assign out[89] = in[350];
    assign out[287] = in[351];
    assign out[138] = in[352];
    assign out[579] = in[353];
    assign out[206] = in[354];
    assign out[271] = in[355];
    assign out[142] = in[356];
    assign out[179] = in[357];
    assign out[274] = in[358];
    assign out[145] = in[359];
    assign out[390] = in[360];
    assign out[621] = in[361];
    assign out[248] = in[362];
    assign out[52] = in[363];
    assign out[266] = in[364];
    assign out[291] = in[365];
    assign out[366] = in[366];
    assign out[573] = in[367];
    assign out[563] = in[368];
    assign out[58] = in[369];
    assign out[17] = in[370];
    assign out[183] = in[371];
    assign out[111] = in[372];
    assign out[225] = in[373];
    assign out[403] = in[374];
    assign out[340] = in[375];
    assign out[1] = in[376];
    assign out[627] = in[377];
    assign out[396] = in[378];
    assign out[118] = in[379];
    assign out[512] = in[380];
    assign out[2] = in[381];
    assign out[413] = in[382];
    assign out[275] = in[383];
    assign out[587] = in[384];
    assign out[483] = in[385];
    assign out[346] = in[386];
    assign out[85] = in[387];
    assign out[198] = in[388];
    assign out[63] = in[389];
    assign out[219] = in[390];
    assign out[268] = in[391];
    assign out[427] = in[392];
    assign out[534] = in[393];
    assign out[114] = in[394];
    assign out[160] = in[395];
    assign out[149] = in[396];
    assign out[433] = in[397];
    assign out[294] = in[398];
    assign out[424] = in[399];
    assign out[547] = in[400];
    assign out[361] = in[401];
    assign out[82] = in[402];
    assign out[95] = in[403];
    assign out[503] = in[404];
    assign out[326] = in[405];
    assign out[13] = in[406];
    assign out[469] = in[407];
    assign out[620] = in[408];
    assign out[342] = in[409];
    assign out[625] = in[410];
    assign out[449] = in[411];
    assign out[603] = in[412];
    assign out[84] = in[413];
    assign out[450] = in[414];
    assign out[180] = in[415];
    assign out[233] = in[416];
    assign out[190] = in[417];
    assign out[261] = in[418];
    assign out[457] = in[419];
    assign out[166] = in[420];
    assign out[560] = in[421];
    assign out[93] = in[422];
    assign out[638] = in[423];
    assign out[237] = in[424];
    assign out[123] = in[425];
    assign out[199] = in[426];
    assign out[463] = in[427];
    assign out[20] = in[428];
    assign out[570] = in[429];
    assign out[402] = in[430];
    assign out[59] = in[431];
    assign out[133] = in[432];
    assign out[302] = in[433];
    assign out[375] = in[434];
    assign out[27] = in[435];
    assign out[513] = in[436];
    assign out[306] = in[437];
    assign out[68] = in[438];
    assign out[110] = in[439];
    assign out[515] = in[440];
    assign out[608] = in[441];
    assign out[338] = in[442];
    assign out[50] = in[443];
    assign out[10] = in[444];
    assign out[61] = in[445];
    assign out[471] = in[446];
    assign out[316] = in[447];
    assign out[317] = in[448];
    assign out[511] = in[449];
    assign out[16] = in[450];
    assign out[216] = in[451];
    assign out[141] = in[452];
    assign out[258] = in[453];
    assign out[286] = in[454];
    assign out[7] = in[455];
    assign out[112] = in[456];
    assign out[67] = in[457];
    assign out[88] = in[458];
    assign out[51] = in[459];
    assign out[599] = in[460];
    assign out[357] = in[461];
    assign out[26] = in[462];
    assign out[370] = in[463];
    assign out[74] = in[464];
    assign out[230] = in[465];
    assign out[550] = in[466];
    assign out[594] = in[467];
    assign out[619] = in[468];
    assign out[242] = in[469];
    assign out[223] = in[470];
    assign out[441] = in[471];
    assign out[329] = in[472];
    assign out[330] = in[473];
    assign out[551] = in[474];
    assign out[446] = in[475];
    assign out[559] = in[476];
    assign out[69] = in[477];
    assign out[439] = in[478];
    assign out[336] = in[479];
    assign out[245] = in[480];
    assign out[556] = in[481];
    assign out[378] = in[482];
    assign out[455] = in[483];
    assign out[30] = in[484];
    assign out[612] = in[485];
    assign out[589] = in[486];
    assign out[634] = in[487];
    assign out[636] = in[488];
    assign out[358] = in[489];
    assign out[120] = in[490];
    assign out[200] = in[491];
    assign out[567] = in[492];
    assign out[532] = in[493];
    assign out[243] = in[494];
    assign out[65] = in[495];
    assign out[623] = in[496];
    assign out[581] = in[497];
    assign out[143] = in[498];
    assign out[376] = in[499];
    assign out[28] = in[500];
    assign out[398] = in[501];
    assign out[334] = in[502];
    assign out[188] = in[503];
    assign out[543] = in[504];
    assign out[516] = in[505];
    assign out[590] = in[506];
    assign out[53] = in[507];
    assign out[36] = in[508];
    assign out[146] = in[509];
    assign out[76] = in[510];
    assign out[132] = in[511];
    assign out[195] = in[512];
    assign out[152] = in[513];
    assign out[289] = in[514];
    assign out[15] = in[515];
    assign out[437] = in[516];
    assign out[136] = in[517];
    assign out[305] = in[518];
    assign out[473] = in[519];
    assign out[381] = in[520];
    assign out[192] = in[521];
    assign out[161] = in[522];
    assign out[374] = in[523];
    assign out[509] = in[524];
    assign out[73] = in[525];
    assign out[301] = in[526];
    assign out[150] = in[527];
    assign out[419] = in[528];
    assign out[401] = in[529];
    assign out[420] = in[530];
    assign out[259] = in[531];
    assign out[126] = in[532];
    assign out[578] = in[533];
    assign out[18] = in[534];
    assign out[278] = in[535];
    assign out[408] = in[536];
    assign out[492] = in[537];
    assign out[22] = in[538];
    assign out[87] = in[539];
    assign out[211] = in[540];
    assign out[212] = in[541];
    assign out[8] = in[542];
    assign out[391] = in[543];
    assign out[307] = in[544];
    assign out[238] = in[545];
    assign out[478] = in[546];
    assign out[47] = in[547];
    assign out[94] = in[548];
    assign out[311] = in[549];
    assign out[486] = in[550];
    assign out[33] = in[551];
    assign out[464] = in[552];
    assign out[128] = in[553];
    assign out[159] = in[554];
    assign out[130] = in[555];
    assign out[86] = in[556];
    assign out[602] = in[557];
    assign out[385] = in[558];
    assign out[282] = in[559];
    assign out[386] = in[560];
    assign out[107] = in[561];
    assign out[92] = in[562];
    assign out[524] = in[563];
    assign out[392] = in[564];
    assign out[194] = in[565];
    assign out[205] = in[566];
    assign out[97] = in[567];
    assign out[98] = in[568];
    assign out[5] = in[569];
    assign out[253] = in[570];
    assign out[119] = in[571];
    assign out[283] = in[572];
    assign out[148] = in[573];
    assign out[285] = in[574];
    assign out[140] = in[575];
    assign out[617] = in[576];
    assign out[558] = in[577];
    assign out[575] = in[578];
    assign out[109] = in[579];
    assign out[377] = in[580];
    assign out[626] = in[581];
    assign out[607] = in[582];
    assign out[113] = in[583];
    assign out[4] = in[584];
    assign out[372] = in[585];
    assign out[454] = in[586];
    assign out[568] = in[587];
    assign out[217] = in[588];
    assign out[164] = in[589];
    assign out[229] = in[590];
    assign out[9] = in[591];
    assign out[197] = in[592];
    assign out[232] = in[593];
    assign out[387] = in[594];
    assign out[528] = in[595];
    assign out[529] = in[596];
    assign out[425] = in[597];
    assign out[537] = in[598];
    assign out[491] = in[599];
    assign out[299] = in[600];
    assign out[409] = in[601];
    assign out[428] = in[602];
    assign out[493] = in[603];
    assign out[273] = in[604];
    assign out[495] = in[605];
    assign out[368] = in[606];
    assign out[276] = in[607];
    assign out[272] = in[608];
    assign out[320] = in[609];
    assign out[436] = in[610];
    assign out[415] = in[611];
    assign out[96] = in[612];
    assign out[79] = in[613];
    assign out[505] = in[614];
    assign out[158] = in[615];
    assign out[549] = in[616];
    assign out[465] = in[617];
    assign out[129] = in[618];
    assign out[580] = in[619];
    assign out[384] = in[620];
    assign out[290] = in[621];
    assign out[163] = in[622];
    assign out[246] = in[623];
    assign out[44] = in[624];
    assign out[353] = in[625];
    assign out[255] = in[626];
    assign out[630] = in[627];
    assign out[169] = in[628];
    assign out[610] = in[629];
    assign out[277] = in[630];
    assign out[250] = in[631];
    assign out[331] = in[632];
    assign out[176] = in[633];
    assign out[100] = in[634];
    assign out[564] = in[635];
    assign out[359] = in[636];
    assign out[380] = in[637];
    assign out[371] = in[638];
    assign out[536] = in[639];
endmodule

module odo_apply_pbox1(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[6] = in[0];
    assign out[484] = in[1];
    assign out[367] = in[2];
    assign out[347] = in[3];
    assign out[69] = in[4];
    assign out[597] = in[5];
    assign out[68] = in[6];
    assign out[112] = in[7];
    assign out[73] = in[8];
    assign out[380] = in[9];
    assign out[429] = in[10];
    assign out[508] = in[11];
    assign out[140] = in[12];
    assign out[296] = in[13];
    assign out[617] = in[14];
    assign out[458] = in[15];
    assign out[385] = in[16];
    assign out[130] = in[17];
    assign out[384] = in[18];
    assign out[547] = in[19];
    assign out[613] = in[20];
    assign out[185] = in[21];
    assign out[604] = in[22];
    assign out[266] = in[23];
    assign out[467] = in[24];
    assign out[2] = in[25];
    assign out[57] = in[26];
    assign out[4] = in[27];
    assign out[407] = in[28];
    assign out[99] = in[29];
    assign out[193] = in[30];
    assign out[144] = in[31];
    assign out[550] = in[32];
    assign out[31] = in[33];
    assign out[104] = in[34];
    assign out[33] = in[35];
    assign out[565] = in[36];
    assign out[280] = in[37];
    assign out[526] = in[38];
    assign out[340] = in[39];
    assign out[343] = in[40];
    assign out[486] = in[41];
    assign out[43] = in[42];
    assign out[235] = in[43];
    assign out[324] = in[44];
    assign out[348] = in[45];
    assign out[283] = in[46];
    assign out[466] = in[47];
    assign out[417] = in[48];
    assign out[428] = in[49];
    assign out[238] = in[50];
    assign out[164] = in[51];
    assign out[631] = in[52];
    assign out[54] = in[53];
    assign out[153] = in[54];
    assign out[410] = in[55];
    assign out[638] = in[56];
    assign out[24] = in[57];
    assign out[113] = in[58];
    assign out[302] = in[59];
    assign out[361] = in[60];
    assign out[28] = in[61];
    assign out[29] = in[62];
    assign out[247] = in[63];
    assign out[445] = in[64];
    assign out[56] = in[65];
    assign out[485] = in[66];
    assign out[446] = in[67];
    assign out[498] = in[68];
    assign out[488] = in[69];
    assign out[371] = in[70];
    assign out[308] = in[71];
    assign out[600] = in[72];
    assign out[255] = in[73];
    assign out[602] = in[74];
    assign out[494] = in[75];
    assign out[530] = in[76];
    assign out[394] = in[77];
    assign out[529] = in[78];
    assign out[199] = in[79];
    assign out[204] = in[80];
    assign out[260] = in[81];
    assign out[533] = in[82];
    assign out[262] = in[83];
    assign out[125] = in[84];
    assign out[83] = in[85];
    assign out[401] = in[86];
    assign out[64] = in[87];
    assign out[542] = in[88];
    assign out[513] = in[89];
    assign out[3] = in[90];
    assign out[190] = in[91];
    assign out[473] = in[92];
    assign out[448] = in[93];
    assign out[409] = in[94];
    assign out[155] = in[95];
    assign out[475] = in[96];
    assign out[561] = in[97];
    assign out[197] = in[98];
    assign out[628] = in[99];
    assign out[551] = in[100];
    assign out[320] = in[101];
    assign out[326] = in[102];
    assign out[420] = in[103];
    assign out[46] = in[104];
    assign out[82] = in[105];
    assign out[142] = in[106];
    assign out[108] = in[107];
    assign out[236] = in[108];
    assign out[333] = in[109];
    assign out[44] = in[110];
    assign out[160] = in[111];
    assign out[470] = in[112];
    assign out[114] = in[113];
    assign out[287] = in[114];
    assign out[432] = in[115];
    assign out[107] = in[116];
    assign out[171] = in[117];
    assign out[154] = in[118];
    assign out[168] = in[119];
    assign out[344] = in[120];
    assign out[358] = in[121];
    assign out[221] = in[122];
    assign out[36] = in[123];
    assign out[58] = in[124];
    assign out[440] = in[125];
    assign out[492] = in[126];
    assign out[591] = in[127];
    assign out[227] = in[128];
    assign out[393] = in[129];
    assign out[129] = in[130];
    assign out[161] = in[131];
    assign out[345] = in[132];
    assign out[584] = in[133];
    assign out[517] = in[134];
    assign out[399] = in[135];
    assign out[523] = in[136];
    assign out[489] = in[137];
    assign out[522] = in[138];
    assign out[559] = in[139];
    assign out[605] = in[140];
    assign out[323] = in[141];
    assign out[120] = in[142];
    assign out[594] = in[143];
    assign out[609] = in[144];
    assign out[241] = in[145];
    assign out[49] = in[146];
    assign out[400] = in[147];
    assign out[126] = in[148];
    assign out[285] = in[149];
    assign out[570] = in[150];
    assign out[538] = in[151];
    assign out[603] = in[152];
    assign out[537] = in[153];
    assign out[354] = in[154];
    assign out[65] = in[155];
    assign out[305] = in[156];
    assign out[474] = in[157];
    assign out[500] = in[158];
    assign out[546] = in[159];
    assign out[200] = in[160];
    assign out[544] = in[161];
    assign out[311] = in[162];
    assign out[17] = in[163];
    assign out[481] = in[164];
    assign out[184] = in[165];
    assign out[80] = in[166];
    assign out[303] = in[167];
    assign out[555] = in[168];
    assign out[18] = in[169];
    assign out[624] = in[170];
    assign out[201] = in[171];
    assign out[637] = in[172];
    assign out[464] = in[173];
    assign out[209] = in[174];
    assign out[141] = in[175];
    assign out[378] = in[176];
    assign out[437] = in[177];
    assign out[438] = in[178];
    assign out[535] = in[179];
    assign out[220] = in[180];
    assign out[136] = in[181];
    assign out[636] = in[182];
    assign out[365] = in[183];
    assign out[472] = in[184];
    assign out[449] = in[185];
    assign out[587] = in[186];
    assign out[574] = in[187];
    assign out[363] = in[188];
    assign out[480] = in[189];
    assign out[450] = in[190];
    assign out[592] = in[191];
    assign out[639] = in[192];
    assign out[169] = in[193];
    assign out[520] = in[194];
    assign out[150] = in[195];
    assign out[579] = in[196];
    assign out[580] = in[197];
    assign out[47] = in[198];
    assign out[589] = in[199];
    assign out[583] = in[200];
    assign out[273] = in[201];
    assign out[416] = in[202];
    assign out[42] = in[203];
    assign out[418] = in[204];
    assign out[496] = in[205];
    assign out[355] = in[206];
    assign out[117] = in[207];
    assign out[499] = in[208];
    assign out[249] = in[209];
    assign out[593] = in[210];
    assign out[121] = in[211];
    assign out[426] = in[212];
    assign out[232] = in[213];
    assign out[63] = in[214];
    assign out[598] = in[215];
    assign out[290] = in[216];
    assign out[540] = in[217];
    assign out[173] = in[218];
    assign out[330] = in[219];
    assign out[539] = in[220];
    assign out[295] = in[221];
    assign out[482] = in[222];
    assign out[191] = in[223];
    assign out[282] = in[224];
    assign out[548] = in[225];
    assign out[364] = in[226];
    assign out[519] = in[227];
    assign out[286] = in[228];
    assign out[276] = in[229];
    assign out[366] = in[230];
    assign out[77] = in[231];
    assign out[633] = in[232];
    assign out[457] = in[233];
    assign out[288] = in[234];
    assign out[139] = in[235];
    assign out[425] = in[236];
    assign out[497] = in[237];
    assign out[502] = in[238];
    assign out[207] = in[239];
    assign out[312] = in[240];
    assign out[352] = in[241];
    assign out[91] = in[242];
    assign out[379] = in[243];
    assign out[243] = in[244];
    assign out[211] = in[245];
    assign out[32] = in[246];
    assign out[332] = in[247];
    assign out[462] = in[248];
    assign out[270] = in[249];
    assign out[413] = in[250];
    assign out[219] = in[251];
    assign out[388] = in[252];
    assign out[545] = in[253];
    assign out[225] = in[254];
    assign out[405] = in[255];
    assign out[179] = in[256];
    assign out[230] = in[257];
    assign out[532] = in[258];
    assign out[127] = in[259];
    assign out[251] = in[260];
    assign out[325] = in[261];
    assign out[189] = in[262];
    assign out[611] = in[263];
    assign out[186] = in[264];
    assign out[252] = in[265];
    assign out[614] = in[266];
    assign out[477] = in[267];
    assign out[493] = in[268];
    assign out[119] = in[269];
    assign out[192] = in[270];
    assign out[618] = in[271];
    assign out[291] = in[272];
    assign out[131] = in[273];
    assign out[629] = in[274];
    assign out[76] = in[275];
    assign out[373] = in[276];
    assign out[341] = in[277];
    assign out[375] = in[278];
    assign out[19] = in[279];
    assign out[143] = in[280];
    assign out[208] = in[281];
    assign out[406] = in[282];
    assign out[521] = in[283];
    assign out[165] = in[284];
    assign out[377] = in[285];
    assign out[23] = in[286];
    assign out[315] = in[287];
    assign out[571] = in[288];
    assign out[216] = in[289];
    assign out[105] = in[290];
    assign out[501] = in[291];
    assign out[215] = in[292];
    assign out[93] = in[293];
    assign out[567] = in[294];
    assign out[632] = in[295];
    assign out[278] = in[296];
    assign out[588] = in[297];
    assign out[444] = in[298];
    assign out[573] = in[299];
    assign out[145] = in[300];
    assign out[87] = in[301];
    assign out[585] = in[302];
    assign out[118] = in[303];
    assign out[304] = in[304];
    assign out[543] = in[305];
    assign out[608] = in[306];
    assign out[495] = in[307];
    assign out[40] = in[308];
    assign out[182] = in[309];
    assign out[356] = in[310];
    assign out[453] = in[311];
    assign out[157] = in[312];
    assign out[424] = in[313];
    assign out[187] = in[314];
    assign out[51] = in[315];
    assign out[256] = in[316];
    assign out[226] = in[317];
    assign out[5] = in[318];
    assign out[461] = in[319];
    assign out[7] = in[320];
    assign out[612] = in[321];
    assign out[549] = in[322];
    assign out[59] = in[323];
    assign out[626] = in[324];
    assign out[439] = in[325];
    assign out[536] = in[326];
    assign out[610] = in[327];
    assign out[374] = in[328];
    assign out[202] = in[329];
    assign out[67] = in[330];
    assign out[541] = in[331];
    assign out[507] = in[332];
    assign out[430] = in[333];
    assign out[338] = in[334];
    assign out[86] = in[335];
    assign out[135] = in[336];
    assign out[196] = in[337];
    assign out[307] = in[338];
    assign out[386] = in[339];
    assign out[203] = in[340];
    assign out[250] = in[341];
    assign out[516] = in[342];
    assign out[1] = in[343];
    assign out[518] = in[344];
    assign out[564] = in[345];
    assign out[346] = in[346];
    assign out[205] = in[347];
    assign out[84] = in[348];
    assign out[576] = in[349];
    assign out[319] = in[350];
    assign out[578] = in[351];
    assign out[321] = in[352];
    assign out[562] = in[353];
    assign out[217] = in[354];
    assign out[337] = in[355];
    assign out[229] = in[356];
    assign out[293] = in[357];
    assign out[34] = in[358];
    assign out[27] = in[359];
    assign out[300] = in[360];
    assign out[224] = in[361];
    assign out[98] = in[362];
    assign out[95] = in[363];
    assign out[163] = in[364];
    assign out[369] = in[365];
    assign out[490] = in[366];
    assign out[322] = in[367];
    assign out[149] = in[368];
    assign out[515] = in[369];
    assign out[590] = in[370];
    assign out[389] = in[371];
    assign out[166] = in[372];
    assign out[172] = in[373];
    assign out[471] = in[374];
    assign out[97] = in[375];
    assign out[239] = in[376];
    assign out[268] = in[377];
    assign out[237] = in[378];
    assign out[178] = in[379];
    assign out[38] = in[380];
    assign out[272] = in[381];
    assign out[55] = in[382];
    assign out[228] = in[383];
    assign out[625] = in[384];
    assign out[188] = in[385];
    assign out[147] = in[386];
    assign out[12] = in[387];
    assign out[505] = in[388];
    assign out[566] = in[389];
    assign out[621] = in[390];
    assign out[101] = in[391];
    assign out[569] = in[392];
    assign out[218] = in[393];
    assign out[524] = in[394];
    assign out[20] = in[395];
    assign out[382] = in[396];
    assign out[478] = in[397];
    assign out[11] = in[398];
    assign out[257] = in[399];
    assign out[110] = in[400];
    assign out[514] = in[401];
    assign out[455] = in[402];
    assign out[318] = in[403];
    assign out[132] = in[404];
    assign out[21] = in[405];
    assign out[45] = in[406];
    assign out[601] = in[407];
    assign out[404] = in[408];
    assign out[510] = in[409];
    assign out[586] = in[410];
    assign out[88] = in[411];
    assign out[89] = in[412];
    assign out[148] = in[413];
    assign out[213] = in[414];
    assign out[240] = in[415];
    assign out[469] = in[416];
    assign out[328] = in[417];
    assign out[615] = in[418];
    assign out[158] = in[419];
    assign out[267] = in[420];
    assign out[534] = in[421];
    assign out[269] = in[422];
    assign out[572] = in[423];
    assign out[223] = in[424];
    assign out[41] = in[425];
    assign out[284] = in[426];
    assign out[70] = in[427];
    assign out[398] = in[428];
    assign out[463] = in[429];
    assign out[281] = in[430];
    assign out[607] = in[431];
    assign out[231] = in[432];
    assign out[563] = in[433];
    assign out[90] = in[434];
    assign out[81] = in[435];
    assign out[331] = in[436];
    assign out[134] = in[437];
    assign out[292] = in[438];
    assign out[174] = in[439];
    assign out[362] = in[440];
    assign out[554] = in[441];
    assign out[122] = in[442];
    assign out[242] = in[443];
    assign out[100] = in[444];
    assign out[575] = in[445];
    assign out[483] = in[446];
    assign out[342] = in[447];
    assign out[94] = in[448];
    assign out[210] = in[449];
    assign out[423] = in[450];
    assign out[309] = in[451];
    assign out[306] = in[452];
    assign out[35] = in[453];
    assign out[15] = in[454];
    assign out[183] = in[455];
    assign out[8] = in[456];
    assign out[103] = in[457];
    assign out[451] = in[458];
    assign out[381] = in[459];
    assign out[263] = in[460];
    assign out[13] = in[461];
    assign out[37] = in[462];
    assign out[314] = in[463];
    assign out[212] = in[464];
    assign out[397] = in[465];
    assign out[244] = in[466];
    assign out[298] = in[467];
    assign out[60] = in[468];
    assign out[133] = in[469];
    assign out[248] = in[470];
    assign out[206] = in[471];
    assign out[115] = in[472];
    assign out[116] = in[473];
    assign out[264] = in[474];
    assign out[50] = in[475];
    assign out[279] = in[476];
    assign out[52] = in[477];
    assign out[265] = in[478];
    assign out[310] = in[479];
    assign out[334] = in[480];
    assign out[30] = in[481];
    assign out[411] = in[482];
    assign out[350] = in[483];
    assign out[390] = in[484];
    assign out[316] = in[485];
    assign out[78] = in[486];
    assign out[277] = in[487];
    assign out[335] = in[488];
    assign out[619] = in[489];
    assign out[479] = in[490];
    assign out[557] = in[491];
    assign out[622] = in[492];
    assign out[606] = in[493];
    assign out[261] = in[494];
    assign out[427] = in[495];
    assign out[75] = in[496];
    assign out[630] = in[497];
    assign out[246] = in[498];
    assign out[74] = in[499];
    assign out[351] = in[500];
    assign out[53] = in[501];
    assign out[431] = in[502];
    assign out[392] = in[503];
    assign out[525] = in[504];
    assign out[180] = in[505];
    assign out[435] = in[506];
    assign out[396] = in[507];
    assign out[128] = in[508];
    assign out[376] = in[509];
    assign out[25] = in[510];
    assign out[436] = in[511];
    assign out[422] = in[512];
    assign out[123] = in[513];
    assign out[558] = in[514];
    assign out[476] = in[515];
    assign out[175] = in[516];
    assign out[349] = in[517];
    assign out[454] = in[518];
    assign out[62] = in[519];
    assign out[468] = in[520];
    assign out[0] = in[521];
    assign out[124] = in[522];
    assign out[329] = in[523];
    assign out[568] = in[524];
    assign out[531] = in[525];
    assign out[48] = in[526];
    assign out[176] = in[527];
    assign out[289] = in[528];
    assign out[465] = in[529];
    assign out[336] = in[530];
    assign out[620] = in[531];
    assign out[274] = in[532];
    assign out[156] = in[533];
    assign out[66] = in[534];
    assign out[253] = in[535];
    assign out[9] = in[536];
    assign out[447] = in[537];
    assign out[357] = in[538];
    assign out[61] = in[539];
    assign out[22] = in[540];
    assign out[146] = in[541];
    assign out[85] = in[542];
    assign out[491] = in[543];
    assign out[553] = in[544];
    assign out[433] = in[545];
    assign out[151] = in[546];
    assign out[353] = in[547];
    assign out[528] = in[548];
    assign out[198] = in[549];
    assign out[511] = in[550];
    assign out[275] = in[551];
    assign out[10] = in[552];
    assign out[138] = in[553];
    assign out[560] = in[554];
    assign out[301] = in[555];
    assign out[317] = in[556];
    assign out[222] = in[557];
    assign out[245] = in[558];
    assign out[102] = in[559];
    assign out[39] = in[560];
    assign out[634] = in[561];
    assign out[259] = in[562];
    assign out[460] = in[563];
    assign out[233] = in[564];
    assign out[635] = in[565];
    assign out[599] = in[566];
    assign out[254] = in[567];
    assign out[26] = in[568];
    assign out[106] = in[569];
    assign out[595] = in[570];
    assign out[577] = in[571];
    assign out[195] = in[572];
    assign out[111] = in[573];
    assign out[271] = in[574];
    assign out[459] = in[575];
    assign out[556] = in[576];
    assign out[487] = in[577];
    assign out[372] = in[578];
    assign out[403] = in[579];
    assign out[258] = in[580];
    assign out[327] = in[581];
    assign out[370] = in[582];
    assign out[313] = in[583];
    assign out[339] = in[584];
    assign out[527] = in[585];
    assign out[181] = in[586];
    assign out[395] = in[587];
    assign out[421] = in[588];
    assign out[71] = in[589];
    assign out[414] = in[590];
    assign out[616] = in[591];
    assign out[177] = in[592];
    assign out[72] = in[593];
    assign out[402] = in[594];
    assign out[299] = in[595];
    assign out[442] = in[596];
    assign out[443] = in[597];
    assign out[623] = in[598];
    assign out[360] = in[599];
    assign out[503] = in[600];
    assign out[581] = in[601];
    assign out[441] = in[602];
    assign out[506] = in[603];
    assign out[359] = in[604];
    assign out[387] = in[605];
    assign out[137] = in[606];
    assign out[415] = in[607];
    assign out[167] = in[608];
    assign out[194] = in[609];
    assign out[552] = in[610];
    assign out[79] = in[611];
    assign out[16] = in[612];
    assign out[582] = in[613];
    assign out[434] = in[614];
    assign out[383] = in[615];
    assign out[504] = in[616];
    assign out[96] = in[617];
    assign out[159] = in[618];
    assign out[92] = in[619];
    assign out[14] = in[620];
    assign out[627] = in[621];
    assign out[391] = in[622];
    assign out[456] = in[623];
    assign out[214] = in[624];
    assign out[509] = in[625];
    assign out[152] = in[626];
    assign out[596] = in[627];
    assign out[294] = in[628];
    assign out[170] = in[629];
    assign out[412] = in[630];
    assign out[297] = in[631];
    assign out[452] = in[632];
    assign out[234] = in[633];
    assign out[512] = in[634];
    assign out[109] = in[635];
    assign out[162] = in[636];
    assign out[419] = in[637];
    assign out[368] = in[638];
    assign out[408] = in[639];
endmodule

module odo_rotation_helper(in, out);
    input [63:0] in;
    output [63:0] out;
    assign out = {in[30:0], in[63:31]} ^ {in[39:0], in[63:40]} ^ {in[40:0], in[63:41]} ^ {in[1:0], in[63:2]} ^ {in[21:0], in[63:22]} ^ {in[20:0], in[63:21]};
endmodule

module odo_apply_rotations(in, out);
    input [639:0] in;
    output [639:0] out;
    wire [639:0] rot;
    odo_rotation_helper rot0inst(in[63:0], rot[63:0]);
    odo_rotation_helper rot1inst(in[127:64], rot[127:64]);
    odo_rotation_helper rot2inst(in[191:128], rot[191:128]);
    odo_rotation_helper rot3inst(in[255:192], rot[255:192]);
    odo_rotation_helper rot4inst(in[319:256], rot[319:256]);
    odo_rotation_helper rot5inst(in[383:320], rot[383:320]);
    odo_rotation_helper rot6inst(in[447:384], rot[447:384]);
    odo_rotation_helper rot7inst(in[511:448], rot[511:448]);
    odo_rotation_helper rot8inst(in[575:512], rot[575:512]);
    odo_rotation_helper rot9inst(in[639:576], rot[639:576]);
    assign out = rot ^ {in[63:0], in[639:64]};
endmodule

module odo_apply_round_key(key, in, out);
    input [9:0] key;
    input [639:0] in;
    output [639:0] out;
    assign out[0] = in[0] ^ key[0];
    assign out[63:1] = in[63:1];
    assign out[64] = in[64] ^ key[1];
    assign out[127:65] = in[127:65];
    assign out[128] = in[128] ^ key[2];
    assign out[191:129] = in[191:129];
    assign out[192] = in[192] ^ key[3];
    assign out[255:193] = in[255:193];
    assign out[256] = in[256] ^ key[4];
    assign out[319:257] = in[319:257];
    assign out[320] = in[320] ^ key[5];
    assign out[383:321] = in[383:321];
    assign out[384] = in[384] ^ key[6];
    assign out[447:385] = in[447:385];
    assign out[448] = in[448] ^ key[7];
    assign out[511:449] = in[511:449];
    assign out[512] = in[512] ^ key[8];
    assign out[575:513] = in[575:513];
    assign out[576] = in[576] ^ key[9];
    assign out[639:577] = in[639:577];
endmodule

module odo_full_round(clk, roundkey, in, out);
    input clk;
    input [9:0] roundkey;
    input [639:0] in;
    output [639:0] out;
    wire [639:0] mid[0:3];
    odo_apply_pbox0 pbox0inst(in, mid[0]);
    odo_apply_sboxes sboxes(clk, mid[0], mid[1]);
    odo_apply_pbox1 pbox1inst(mid[1], mid[2]);
    odo_apply_rotations rotations(mid[2], mid[3]);
    odo_apply_round_key keys(roundkey, mid[3], out);
endmodule

module odo_get_round_key0(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h0b5;
        4'h1: key <= 10'h0d3;
        4'h2: key <= 10'h26c;
        4'h3: key <= 10'h1ad;
        4'h4: key <= 10'h360;
        4'h5: key <= 10'h2d4;
        4'h6: key <= 10'h2b2;
        4'h7: key <= 10'h287;
        4'h8: key <= 10'h24f;
        4'h9: key <= 10'h360;
    endcase
    end
endmodule

module odo_get_round_key1(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h10e;
        4'h1: key <= 10'h0c1;
        4'h2: key <= 10'h120;
        4'h3: key <= 10'h21d;
        4'h4: key <= 10'h311;
        4'h5: key <= 10'h240;
        4'h6: key <= 10'h366;
        4'h7: key <= 10'h3c6;
        4'h8: key <= 10'h2e2;
        4'h9: key <= 10'h144;
    endcase
    end
endmodule

module odo_get_round_key2(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h3ef;
        4'h1: key <= 10'h2d9;
        4'h2: key <= 10'h2d7;
        4'h3: key <= 10'h229;
        4'h4: key <= 10'h008;
        4'h5: key <= 10'h335;
        4'h6: key <= 10'h091;
        4'h7: key <= 10'h073;
        4'h8: key <= 10'h1ce;
        4'h9: key <= 10'h1c6;
    endcase
    end
endmodule

module odo_get_round_key3(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h02b;
        4'h1: key <= 10'h1e1;
        4'h2: key <= 10'h340;
        4'h3: key <= 10'h3c7;
        4'h4: key <= 10'h0a6;
        4'h5: key <= 10'h0b2;
        4'h6: key <= 10'h223;
        4'h7: key <= 10'h2fb;
        4'h8: key <= 10'h3d7;
    endcase
    end
endmodule

module odo_get_round_key4(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h2d1;
        4'h1: key <= 10'h081;
        4'h2: key <= 10'h0fd;
        4'h3: key <= 10'h080;
        4'h4: key <= 10'h1c4;
        4'h5: key <= 10'h1d6;
        4'h6: key <= 10'h2cf;
        4'h7: key <= 10'h25d;
        4'h8: key <= 10'h083;
    endcase
    end
endmodule

module odo_get_round_key5(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h343;
        4'h1: key <= 10'h227;
        4'h2: key <= 10'h033;
        4'h3: key <= 10'h3ec;
        4'h4: key <= 10'h07b;
        4'h5: key <= 10'h357;
        4'h6: key <= 10'h18c;
        4'h7: key <= 10'h1d6;
        4'h8: key <= 10'h046;
    endcase
    end
endmodule

module odo_get_round_key6(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h2f8;
        4'h1: key <= 10'h290;
        4'h2: key <= 10'h2cb;
        4'h3: key <= 10'h14c;
        4'h4: key <= 10'h185;
        4'h5: key <= 10'h3c2;
        4'h6: key <= 10'h1ab;
        4'h7: key <= 10'h114;
        4'h8: key <= 10'h10d;
    endcase
    end
endmodule

module odo_get_round_key7(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h03b;
        4'h1: key <= 10'h183;
        4'h2: key <= 10'h2cf;
        4'h3: key <= 10'h2dc;
        4'h4: key <= 10'h246;
        4'h5: key <= 10'h0b7;
        4'h6: key <= 10'h1d8;
        4'h7: key <= 10'h2ce;
        4'h8: key <= 10'h3f2;
    endcase
    end
endmodule

module odo_get_round_key8(clk, period, key);
    input clk;
    input [3:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        4'h0: key <= 10'h337;
        4'h1: key <= 10'h36e;
        4'h2: key <= 10'h2ab;
        4'h3: key <= 10'h312;
        4'h4: key <= 10'h312;
        4'h5: key <= 10'h010;
        4'h6: key <= 10'h150;
        4'h7: key <= 10'h0a7;
        4'h8: key <= 10'h0c0;
    endcase
    end
endmodule

module odo_encrypt_loop(clk, in, read, out, write);
    input clk;
    input [639:0] in;
    input read;
    output reg [639:0] out;
    output write;
    reg [639:0] state[9:0];
    wire [639:0] next[9:0];
    always @(posedge clk) state[1] <= next[0];
    always @(posedge clk) state[2] <= next[1];
    always @(posedge clk) state[3] <= next[2];
    always @(posedge clk) state[4] <= next[3];
    always @(posedge clk) state[5] <= next[4];
    always @(posedge clk) state[6] <= next[5];
    always @(posedge clk) state[7] <= next[6];
    always @(posedge clk) state[8] <= next[7];
    always @(posedge clk) state[9] <= next[8];
    assign next[9] = state[9];
    wire [9:0] roundkey[8:0];
    reg [3:0] period[18:0];
    always @(posedge clk) period[1] <= period[0];
    always @(posedge clk) period[2] <= period[1];
    always @(posedge clk) period[3] <= period[2];
    always @(posedge clk) period[4] <= period[3];
    always @(posedge clk) period[5] <= period[4];
    always @(posedge clk) period[6] <= period[5];
    always @(posedge clk) period[7] <= period[6];
    always @(posedge clk) period[8] <= period[7];
    always @(posedge clk) period[9] <= period[8];
    always @(posedge clk) period[10] <= period[9];
    always @(posedge clk) period[11] <= period[10];
    always @(posedge clk) period[12] <= period[11];
    always @(posedge clk) period[13] <= period[12];
    always @(posedge clk) period[14] <= period[13];
    always @(posedge clk) period[15] <= period[14];
    always @(posedge clk) period[16] <= period[15];
    always @(posedge clk) period[17] <= period[16];
    always @(posedge clk) period[18] <= period[17];
    odo_get_round_key0 get_key0(clk, period[0], roundkey[0]);
    odo_full_round round0(clk, roundkey[0], state[0], next[0]);
    odo_get_round_key1 get_key1(clk, period[2], roundkey[1]);
    odo_full_round round1(clk, roundkey[1], state[1], next[1]);
    odo_get_round_key2 get_key2(clk, period[4], roundkey[2]);
    odo_full_round round2(clk, roundkey[2], state[2], next[2]);
    odo_get_round_key3 get_key3(clk, period[6], roundkey[3]);
    odo_full_round round3(clk, roundkey[3], state[3], next[3]);
    odo_get_round_key4 get_key4(clk, period[8], roundkey[4]);
    odo_full_round round4(clk, roundkey[4], state[4], next[4]);
    odo_get_round_key5 get_key5(clk, period[10], roundkey[5]);
    odo_full_round round5(clk, roundkey[5], state[5], next[5]);
    odo_get_round_key6 get_key6(clk, period[12], roundkey[6]);
    odo_full_round round6(clk, roundkey[6], state[6], next[6]);
    odo_get_round_key7 get_key7(clk, period[14], roundkey[7]);
    odo_full_round round7(clk, roundkey[7], state[7], next[7]);
    odo_get_round_key8 get_key8(clk, period[16], roundkey[8]);
    odo_full_round round8(clk, roundkey[8], state[8], next[8]);
    always @(posedge clk) begin
        if (read)
        begin
            period[0] <= 0;
            state[0] <= in;
        end
        else
        begin
            period[0] <= period[18]+1;
            state[0] <= next[9];
        end
        out <= next[2];
    end
    reg [177:0] progress;
    initial progress = 178'h0;
    always @(posedge clk) progress[0] <= read;
    always @(posedge clk) progress[1] <= progress[0];
    always @(posedge clk) progress[2] <= progress[1];
    always @(posedge clk) progress[3] <= progress[2];
    always @(posedge clk) progress[4] <= progress[3];
    always @(posedge clk) progress[5] <= progress[4];
    always @(posedge clk) progress[6] <= progress[5];
    always @(posedge clk) progress[7] <= progress[6];
    always @(posedge clk) progress[8] <= progress[7];
    always @(posedge clk) progress[9] <= progress[8];
    always @(posedge clk) progress[10] <= progress[9];
    always @(posedge clk) progress[11] <= progress[10];
    always @(posedge clk) progress[12] <= progress[11];
    always @(posedge clk) progress[13] <= progress[12];
    always @(posedge clk) progress[14] <= progress[13];
    always @(posedge clk) progress[15] <= progress[14];
    always @(posedge clk) progress[16] <= progress[15];
    always @(posedge clk) progress[17] <= progress[16];
    always @(posedge clk) progress[18] <= progress[17];
    always @(posedge clk) progress[19] <= progress[18];
    always @(posedge clk) progress[20] <= progress[19];
    always @(posedge clk) progress[21] <= progress[20];
    always @(posedge clk) progress[22] <= progress[21];
    always @(posedge clk) progress[23] <= progress[22];
    always @(posedge clk) progress[24] <= progress[23];
    always @(posedge clk) progress[25] <= progress[24];
    always @(posedge clk) progress[26] <= progress[25];
    always @(posedge clk) progress[27] <= progress[26];
    always @(posedge clk) progress[28] <= progress[27];
    always @(posedge clk) progress[29] <= progress[28];
    always @(posedge clk) progress[30] <= progress[29];
    always @(posedge clk) progress[31] <= progress[30];
    always @(posedge clk) progress[32] <= progress[31];
    always @(posedge clk) progress[33] <= progress[32];
    always @(posedge clk) progress[34] <= progress[33];
    always @(posedge clk) progress[35] <= progress[34];
    always @(posedge clk) progress[36] <= progress[35];
    always @(posedge clk) progress[37] <= progress[36];
    always @(posedge clk) progress[38] <= progress[37];
    always @(posedge clk) progress[39] <= progress[38];
    always @(posedge clk) progress[40] <= progress[39];
    always @(posedge clk) progress[41] <= progress[40];
    always @(posedge clk) progress[42] <= progress[41];
    always @(posedge clk) progress[43] <= progress[42];
    always @(posedge clk) progress[44] <= progress[43];
    always @(posedge clk) progress[45] <= progress[44];
    always @(posedge clk) progress[46] <= progress[45];
    always @(posedge clk) progress[47] <= progress[46];
    always @(posedge clk) progress[48] <= progress[47];
    always @(posedge clk) progress[49] <= progress[48];
    always @(posedge clk) progress[50] <= progress[49];
    always @(posedge clk) progress[51] <= progress[50];
    always @(posedge clk) progress[52] <= progress[51];
    always @(posedge clk) progress[53] <= progress[52];
    always @(posedge clk) progress[54] <= progress[53];
    always @(posedge clk) progress[55] <= progress[54];
    always @(posedge clk) progress[56] <= progress[55];
    always @(posedge clk) progress[57] <= progress[56];
    always @(posedge clk) progress[58] <= progress[57];
    always @(posedge clk) progress[59] <= progress[58];
    always @(posedge clk) progress[60] <= progress[59];
    always @(posedge clk) progress[61] <= progress[60];
    always @(posedge clk) progress[62] <= progress[61];
    always @(posedge clk) progress[63] <= progress[62];
    always @(posedge clk) progress[64] <= progress[63];
    always @(posedge clk) progress[65] <= progress[64];
    always @(posedge clk) progress[66] <= progress[65];
    always @(posedge clk) progress[67] <= progress[66];
    always @(posedge clk) progress[68] <= progress[67];
    always @(posedge clk) progress[69] <= progress[68];
    always @(posedge clk) progress[70] <= progress[69];
    always @(posedge clk) progress[71] <= progress[70];
    always @(posedge clk) progress[72] <= progress[71];
    always @(posedge clk) progress[73] <= progress[72];
    always @(posedge clk) progress[74] <= progress[73];
    always @(posedge clk) progress[75] <= progress[74];
    always @(posedge clk) progress[76] <= progress[75];
    always @(posedge clk) progress[77] <= progress[76];
    always @(posedge clk) progress[78] <= progress[77];
    always @(posedge clk) progress[79] <= progress[78];
    always @(posedge clk) progress[80] <= progress[79];
    always @(posedge clk) progress[81] <= progress[80];
    always @(posedge clk) progress[82] <= progress[81];
    always @(posedge clk) progress[83] <= progress[82];
    always @(posedge clk) progress[84] <= progress[83];
    always @(posedge clk) progress[85] <= progress[84];
    always @(posedge clk) progress[86] <= progress[85];
    always @(posedge clk) progress[87] <= progress[86];
    always @(posedge clk) progress[88] <= progress[87];
    always @(posedge clk) progress[89] <= progress[88];
    always @(posedge clk) progress[90] <= progress[89];
    always @(posedge clk) progress[91] <= progress[90];
    always @(posedge clk) progress[92] <= progress[91];
    always @(posedge clk) progress[93] <= progress[92];
    always @(posedge clk) progress[94] <= progress[93];
    always @(posedge clk) progress[95] <= progress[94];
    always @(posedge clk) progress[96] <= progress[95];
    always @(posedge clk) progress[97] <= progress[96];
    always @(posedge clk) progress[98] <= progress[97];
    always @(posedge clk) progress[99] <= progress[98];
    always @(posedge clk) progress[100] <= progress[99];
    always @(posedge clk) progress[101] <= progress[100];
    always @(posedge clk) progress[102] <= progress[101];
    always @(posedge clk) progress[103] <= progress[102];
    always @(posedge clk) progress[104] <= progress[103];
    always @(posedge clk) progress[105] <= progress[104];
    always @(posedge clk) progress[106] <= progress[105];
    always @(posedge clk) progress[107] <= progress[106];
    always @(posedge clk) progress[108] <= progress[107];
    always @(posedge clk) progress[109] <= progress[108];
    always @(posedge clk) progress[110] <= progress[109];
    always @(posedge clk) progress[111] <= progress[110];
    always @(posedge clk) progress[112] <= progress[111];
    always @(posedge clk) progress[113] <= progress[112];
    always @(posedge clk) progress[114] <= progress[113];
    always @(posedge clk) progress[115] <= progress[114];
    always @(posedge clk) progress[116] <= progress[115];
    always @(posedge clk) progress[117] <= progress[116];
    always @(posedge clk) progress[118] <= progress[117];
    always @(posedge clk) progress[119] <= progress[118];
    always @(posedge clk) progress[120] <= progress[119];
    always @(posedge clk) progress[121] <= progress[120];
    always @(posedge clk) progress[122] <= progress[121];
    always @(posedge clk) progress[123] <= progress[122];
    always @(posedge clk) progress[124] <= progress[123];
    always @(posedge clk) progress[125] <= progress[124];
    always @(posedge clk) progress[126] <= progress[125];
    always @(posedge clk) progress[127] <= progress[126];
    always @(posedge clk) progress[128] <= progress[127];
    always @(posedge clk) progress[129] <= progress[128];
    always @(posedge clk) progress[130] <= progress[129];
    always @(posedge clk) progress[131] <= progress[130];
    always @(posedge clk) progress[132] <= progress[131];
    always @(posedge clk) progress[133] <= progress[132];
    always @(posedge clk) progress[134] <= progress[133];
    always @(posedge clk) progress[135] <= progress[134];
    always @(posedge clk) progress[136] <= progress[135];
    always @(posedge clk) progress[137] <= progress[136];
    always @(posedge clk) progress[138] <= progress[137];
    always @(posedge clk) progress[139] <= progress[138];
    always @(posedge clk) progress[140] <= progress[139];
    always @(posedge clk) progress[141] <= progress[140];
    always @(posedge clk) progress[142] <= progress[141];
    always @(posedge clk) progress[143] <= progress[142];
    always @(posedge clk) progress[144] <= progress[143];
    always @(posedge clk) progress[145] <= progress[144];
    always @(posedge clk) progress[146] <= progress[145];
    always @(posedge clk) progress[147] <= progress[146];
    always @(posedge clk) progress[148] <= progress[147];
    always @(posedge clk) progress[149] <= progress[148];
    always @(posedge clk) progress[150] <= progress[149];
    always @(posedge clk) progress[151] <= progress[150];
    always @(posedge clk) progress[152] <= progress[151];
    always @(posedge clk) progress[153] <= progress[152];
    always @(posedge clk) progress[154] <= progress[153];
    always @(posedge clk) progress[155] <= progress[154];
    always @(posedge clk) progress[156] <= progress[155];
    always @(posedge clk) progress[157] <= progress[156];
    always @(posedge clk) progress[158] <= progress[157];
    always @(posedge clk) progress[159] <= progress[158];
    always @(posedge clk) progress[160] <= progress[159];
    always @(posedge clk) progress[161] <= progress[160];
    always @(posedge clk) progress[162] <= progress[161];
    always @(posedge clk) progress[163] <= progress[162];
    always @(posedge clk) progress[164] <= progress[163];
    always @(posedge clk) progress[165] <= progress[164];
    always @(posedge clk) progress[166] <= progress[165];
    always @(posedge clk) progress[167] <= progress[166];
    always @(posedge clk) progress[168] <= progress[167];
    always @(posedge clk) progress[169] <= progress[168];
    always @(posedge clk) progress[170] <= progress[169];
    always @(posedge clk) progress[171] <= progress[170];
    always @(posedge clk) progress[172] <= progress[171];
    always @(posedge clk) progress[173] <= progress[172];
    always @(posedge clk) progress[174] <= progress[173];
    always @(posedge clk) progress[175] <= progress[174];
    always @(posedge clk) progress[176] <= progress[175];
    always @(posedge clk) progress[177] <= progress[176];
    assign write = progress[177];
endmodule

module odo_encrypt(clk, in, read, out, write);
    localparam THROUGHPUT = 10;
    input clk;
    input [639:0] in;
    input read;
    output [639:0] out;
    output write;
    reg [1:0] progress;
    initial progress = 2'h0;
    reg [639:0] state[1:0];
    wire [639:0] next;
    odo_pre_mix premixer(state[0], next);
    odo_encrypt_loop crypter(clk, state[1], progress[1], out, write);
    always @(posedge clk) begin
        progress[0] <= read;
        progress[1] <= progress[0];
        state[0] <= in;
        state[1] <= next;
    end
endmodule
